* netlist generated with vector fitting poles and residues

.subckt total_network node_1 node_2 
X_11 node_1 0 yp11
X_12 node_1 node_2 yp12
X_22 node_2 0 yp22
.ends


* Y'11
.subckt yp11 node_1 0
* Branch 0
Rabr0 node_1 netRa0 414476.48140188813
Lbr0 netRa0 netL0 3.887563647814052e-10
Rbbr0 netL0 0 -1355496.3877445655
Cbr0 netL0 0 7.079979570302878e-22

* Branch 1
Rabr1 node_1 netRa1 595296666.2598804
Lbr1 netRa1 netL1 -7.505893627676451e-09
Rbbr1 netL1 0 -595518367.6129112
Cbr1 netL1 0 -2.1166322460437052e-26

* Branch 2
Rabr2 node_1 netRa2 355756.73483245855
Lbr2 netRa2 netL2 2.580368785481103e-10
Rbbr2 netL2 0 -934716.7388529332
Cbr2 netL2 0 7.893788906612281e-22

* Branch 3
Rabr3 node_1 netRa3 486272.76953370863
Lbr3 netRa3 netL3 2.4394434128439403e-10
Rbbr3 netL3 0 -788614.3834195045
Cbr3 netL3 0 6.434496298243049e-22

* Branch 4
Rabr4 node_1 netRa4 -85257.02826451746
Lbr4 netRa4 netL4 -2.446927895729708e-10
Rbbr4 netL4 0 829155.0676256304
Cbr4 netL4 0 -3.687612325533523e-21

* Branch 5
Rabr5 node_1 netRa5 257809.65565702156
Lbr5 netRa5 netL5 2.3989549430662356e-10
Rbbr5 netL5 0 -980356.916492761
Cbr5 netL5 0 9.67723496347635e-22

* Branch 6
Rabr6 node_1 netRa6 6700707.999203351
Lbr6 netRa6 netL6 -1.401076762238484e-09
Rbbr6 netL6 0 -7322211.643311375
Cbr6 netL6 0 -2.844197618635254e-23

* Branch 7
Rabr7 node_1 netRa7 6714036029.931326
Lbr7 netRa7 netL7 -4.597589538975789e-08
Rbbr7 netL7 0 -6714563511.265519
Cbr7 netL7 0 -1.019705675381903e-27

* Branch 8
Rabr8 node_1 netRa8 4678549.754083234
Lbr8 netRa8 netL8 1.348600847119846e-09
Rbbr8 netL8 0 -5382356.510907061
Cbr8 netL8 0 5.382882402308889e-23

* Branch 9
Rabr9 node_1 netRa9 134217544.16775689
Lbr9 netRa9 netL9 3.503047875847051e-09
Rbbr9 netL9 0 -134480601.83569193
Cbr9 netL9 0 1.9415883752164937e-25

* Branch 10
Rabr10 node_1 netRa10 271420.47237451817
Lbr10 netRa10 netL10 1.777618098689261e-10
Rbbr10 netL10 0 -553478.6912262423
Cbr10 netL10 0 1.1956941020254264e-21

* Branch 11
Rabr11 node_1 netRa11 17449770.1905141
Lbr11 netRa11 netL11 1.1668008456524477e-09
Rbbr11 netL11 0 -17560790.897877827
Cbr11 netL11 0 3.811657479609553e-24

* Branch 12
Rabr12 node_1 netRa12 8968003.159915391
Lbr12 netRa12 netL12 -6.601914246690106e-10
Rbbr12 netL12 0 -9134960.145515803
Cbr12 netL12 0 -8.050007983949907e-24

* Branch 13
Rabr13 node_1 netRa13 6837737.4213986425
Lbr13 netRa13 netL13 9.903356550181433e-10
Rbbr13 netL13 0 -7236441.600988305
Cbr13 netL13 0 2.0056475674949507e-23

* Branch 14
Rabr14 node_1 netRa14 682867.003616919
Lbr14 netRa14 netL14 -4.675057614662034e-10
Rbbr14 netL14 0 -1314629.9591516159
Cbr14 netL14 0 -5.158302415135117e-22

* Branch 15
Rabr15 node_1 netRa15 -1232828.433723843
Lbr15 netRa15 netL15 -6.294261752182286e-10
Rbbr15 netL15 0 1418646.9350645118
Cbr15 netL15 0 -3.619265974398646e-22

* Branch 16
Rabr16 node_1 netRa16 10726826.382466394
Lbr16 netRa16 netL16 1.288741316667207e-09
Rbbr16 netL16 0 -11235642.927088547
Cbr16 netL16 0 1.0706996797645234e-23

* Branch 17
Rabr17 node_1 netRa17 402156.8998362479
Lbr17 netRa17 netL17 -1.930514047272723e-10
Rbbr17 netL17 0 -607108.415142285
Cbr17 netL17 0 -7.865936727840716e-22

* Branch 18
Rabr18 node_1 netRa18 -1354510.3831319248
Lbr18 netRa18 netL18 -6.10398391501598e-10
Rbbr18 netL18 0 1525322.2344613636
Cbr18 netL18 0 -2.9686950091939375e-22

* Branch 19
Rabr19 node_1 netRa19 1620759.6060235214
Lbr19 netRa19 netL19 -5.391790068781643e-10
Rbbr19 netL19 0 -1865032.8359824345
Cbr19 netL19 0 -1.7774754390392288e-22

* Branch 20
Rabr20 node_1 netRa20 3051377.8944083694
Lbr20 netRa20 netL20 -4.672347763098183e-10
Rbbr20 netL20 0 -3164201.938620008
Cbr20 netL20 0 -4.831915036968247e-23

* Branch 21
Rabr21 node_1 netRa21 826624.0794897809
Lbr21 netRa21 netL21 -5.433874631870209e-10
Rbbr21 netL21 0 -1497653.5565640484
Cbr21 netL21 0 -4.361701337028645e-22

* Branch 22
Rabr22 node_1 netRa22 6626.893465684433
Lbr22 netRa22 netL22 1.719903201976538e-10
Rbbr22 netL22 0 -3123020.4442858812
Cbr22 netL22 0 1.0896182664492996e-20

* Branch 23
Rabr23 node_1 netRa23 82602.26149040491
Lbr23 netRa23 netL23 -2.581992685615447e-10
Rbbr23 netL23 0 -582170.7174207667
Cbr23 netL23 0 -5.2243839445175424e-21

* Branch 24
Rabr24 node_1 netRa24 -93140.19931271694
Lbr24 netRa24 netL24 -2.388434942731368e-10
Rbbr24 netL24 0 712047.6002776425
Cbr24 netL24 0 -3.681831975073956e-21

* Branch 25
Rabr25 node_1 netRa25 530451.5031682441
Lbr25 netRa25 netL25 1.499937602595732e-10
Rbbr25 netL25 0 -656652.9552892416
Cbr25 netL25 0 4.316569240409229e-22

* Branch 26
Rabr26 node_1 netRa26 49180.85683124922
Lbr26 netRa26 netL26 3.346442162925014e-11
Rbbr26 netL26 0 -129802.40793730773
Cbr26 netL26 0 5.2723055239519784e-21

* Branch 27
Rabr27 node_1 netRa27 75996.94374488856
Lbr27 netRa27 netL27 1.9843739284380786e-10
Rbbr27 netL27 0 -482807.0830577273
Cbr27 netL27 0 5.51771604225942e-21

* Branch 28
Rabr28 node_1 netRa28 233149.35014725412
Lbr28 netRa28 netL28 -3.5395818812552626e-10
Rbbr28 netL28 0 -601199.6126543933
Cbr28 netL28 0 -2.4974677532651322e-21

* Branch 29
Rabr29 node_1 netRa29 1951701.4963087083
Lbr29 netRa29 netL29 -3.99637014495378e-10
Rbbr29 netL29 0 -2092042.3010939225
Cbr29 netL29 0 -9.773797460847007e-23

* Branch 30
Rabr30 node_1 netRa30 168104.7324078113
Lbr30 netRa30 netL30 -1.9597023489939282e-10
Rbbr30 netL30 0 -523434.14414803113
Cbr30 netL30 0 -2.2104151684316753e-21

* Branch 31
Rabr31 node_1 netRa31 423274.8765852903
Lbr31 netRa31 netL31 1.4842991641871032e-10
Rbbr31 netL31 0 -574973.3563339389
Cbr31 netL31 0 6.11228480254709e-22

* Branch 32
Rabr32 node_1 netRa32 20198164.96034675
Lbr32 netRa32 netL32 -1.1431350696939273e-09
Rbbr32 netL32 0 -20345222.647322938
Cbr32 netL32 0 -2.7808099136193875e-24

* Branch 33
Rabr33 node_1 netRa33 -725244.1963912885
Lbr33 netRa33 netL33 -5.286430833320138e-10
Rbbr33 netL33 0 940144.6871644761
Cbr33 netL33 0 -7.788260043814709e-22

* Branch 34
Rabr34 node_1 netRa34 981378.3297779175
Lbr34 netRa34 netL34 2.1275438071141688e-10
Rbbr34 netL34 0 -1138863.1385261903
Cbr34 netL34 0 1.9060618176400296e-22

* Branch 35
Rabr35 node_1 netRa35 3843936.3132752758
Lbr35 netRa35 netL35 -1.715689073437861e-09
Rbbr35 netL35 0 -5828072.035831923
Cbr35 netL35 0 -7.638367263817796e-23

* Branch 36
Rabr36 node_1 netRa36 2104337.640354159
Lbr36 netRa36 netL36 1.4468533047240664e-09
Rbbr36 netL36 0 -2574475.4894923936
Cbr36 netL36 0 2.6811042997330115e-22

* Branch 37
Rabr37 node_1 netRa37 281663.1725117496
Lbr37 netRa37 netL37 2.62671932859272e-10
Rbbr37 netL37 0 -590652.3755098474
Cbr37 netL37 0 1.5864737765889038e-21

* Branch 38
Rabr38 node_1 netRa38 693220.917856639
Lbr38 netRa38 netL38 -2.124108975368438e-10
Rbbr38 netL38 0 -866608.1403305031
Cbr38 netL38 0 -3.530570550863708e-22

* Branch 39
Rabr39 node_1 netRa39 838779.4211722161
Lbr39 netRa39 netL39 -2.7141582933942407e-10
Rbbr39 netL39 0 -1019539.5611201286
Cbr39 netL39 0 -3.1691081051853113e-22

* Branch 40
Rabr40 node_1 netRa40 884914.2910663267
Lbr40 netRa40 netL40 -2.719662387986462e-10
Rbbr40 netL40 0 -1052874.3708471002
Cbr40 netL40 0 -2.914982381219792e-22

* Branch 41
Rabr41 node_1 netRa41 48068.7688761201
Lbr41 netRa41 netL41 -1.0395892623742593e-10
Rbbr41 netL41 0 -388326.88180937344
Cbr41 netL41 0 -5.515869497025851e-21

* Branch 42
Rabr42 node_1 netRa42 -72253.20469912367
Lbr42 netRa42 netL42 -2.2720507138587039e-10
Rbbr42 netL42 0 798253.295043312
Cbr42 netL42 0 -3.9930573845757844e-21

* Branch 43
Rabr43 node_1 netRa43 921143.2815170797
Lbr43 netRa43 netL43 -2.8700147980718205e-10
Rbbr43 netL43 0 -1091677.638313929
Cbr43 netL43 0 -2.8503120041527567e-22

* Branch 44
Rabr44 node_1 netRa44 2698981.5904697566
Lbr44 netRa44 netL44 8.731625865059637e-10
Rbbr44 netL44 0 -3039090.4857901926
Cbr44 netL44 0 1.0659599832865283e-22

* Branch 45
Rabr45 node_1 netRa45 -218663.70591324675
Lbr45 netRa45 netL45 -2.1475067920314015e-10
Rbbr45 netL45 0 370912.1987428167
Cbr45 netL45 0 -2.6577616868148313e-21

* Branch 46
Rabr46 node_1 netRa46 3392489371.6443124
Lbr46 netRa46 netL46 1.573842684225211e-08
Rbbr46 netL46 0 -3392652445.122111
Cbr46 netL46 0 1.3674481330351707e-27

* Branch 47
Rabr47 node_1 netRa47 -57284.208571625764
Lbr47 netRa47 netL47 2.261534011618886e-10
Rbbr47 netL47 0 654983.0940100783
Cbr47 netL47 0 5.942076237098701e-21

* Branch 48
Rabr48 node_1 netRa48 206798947.48720932
Lbr48 netRa48 netL48 -3.611243459171397e-09
Rbbr48 netL48 0 -206971210.26755908
Cbr48 netL48 0 -8.436712585825185e-26

* Branch 49
Rabr49 node_1 netRa49 -104323.82190539206
Lbr49 netRa49 netL49 -3.921458986533371e-10
Rbbr49 netL49 0 993889.4109562635
Cbr49 netL49 0 -3.825149417514083e-21

* Branch 50
Rabr50 node_1 netRa50 -2111082.1553059714
Lbr50 netRa50 netL50 8.444666921258737e-10
Rbbr50 netL50 0 2285622.9039238296
Cbr50 netL50 0 1.7482861692422948e-22

* Branch 51
Rabr51 node_1 netRa51 -111541.00797511669
Lbr51 netRa51 netL51 -2.26864259411099e-10
Rbbr51 netL51 0 513884.4307375319
Cbr51 netL51 0 -3.978566651125464e-21

* Branch 52
Rabr52 node_1 netRa52 171627.11604617638
Lbr52 netRa52 netL52 1.7199590899612245e-10
Rbbr52 netL52 0 -729080.3871638993
Cbr52 netL52 0 1.3779270587834702e-21

* Branch 53
Rabr53 node_1 netRa53 -632893.307477669
Lbr53 netRa53 netL53 -3.260213032021906e-10
Rbbr53 netL53 0 758577.6106280768
Cbr53 netL53 0 -6.79930762102565e-22

* Branch 54
Rabr54 node_1 netRa54 571944.0408868392
Lbr54 netRa54 netL54 -4.693578841701041e-10
Rbbr54 netL54 0 -1139343.282920003
Cbr54 netL54 0 -7.18983841870224e-22

* Branch 55
Rabr55 node_1 netRa55 1141998.8906765603
Lbr55 netRa55 netL55 -5.594875044329313e-10
Rbbr55 netL55 0 -1587052.8536307472
Cbr55 netL55 0 -3.084205488630102e-22

* Branch 56
Rabr56 node_1 netRa56 837384.5417653923
Lbr56 netRa56 netL56 -3.1277539247756865e-10
Rbbr56 netL56 0 -1142255.2676115595
Cbr56 netL56 0 -3.2677401060605583e-22

* Branch 57
Rabr57 node_1 netRa57 100320257.93287526
Lbr57 netRa57 netL57 -4.331929187582376e-09
Rbbr57 netL57 0 -100650086.95559467
Cbr57 netL57 0 -4.289962081989629e-25

* Branch 58
Rabr58 node_1 netRa58 3989090.994428651
Lbr58 netRa58 netL58 -9.648069305555127e-10
Rbbr58 netL58 0 -4494880.763283733
Cbr58 netL58 0 -5.379151127825912e-23

* Branch 59
Rabr59 node_1 netRa59 203719656.51099873
Lbr59 netRa59 netL59 -6.5615330596806605e-09
Rbbr59 netL59 0 -204166801.78983405
Cbr59 netL59 0 -1.5775050412674639e-25

* Branch 60
Rabr60 node_1 netRa60 4940692.42849858
Lbr60 netRa60 netL60 1.21585083529536e-09
Rbbr60 netL60 0 -5373593.1767965
Cbr60 netL60 0 4.5809176145000313e-23

* Branch 61
Rabr61 node_1 netRa61 7765523.710558203
Lbr61 netRa61 netL61 5.928610949030792e-10
Rbbr61 netL61 0 -7908018.049797745
Cbr61 netL61 0 9.654973618567706e-24

* Branch 62
Rabr62 node_1 netRa62 -583064.3266689259
Lbr62 netRa62 netL62 6.566219132781684e-10
Rbbr62 netL62 0 945879.8649444891
Cbr62 netL62 0 1.189418351700811e-21

* Branch 63
Rabr63 node_1 netRa63 259820.1716123109
Lbr63 netRa63 netL63 4.414549133409172e-10
Rbbr63 netL63 0 -2135272.3592433822
Cbr63 netL63 0 7.9685285654366055e-22

* Branch 64
Rabr64 node_1 netRa64 9041.965634080309
Lbr64 netRa64 netL64 -1.2173828654074592e-10
Rbbr64 netL64 0 -2077425.7860979014
Cbr64 netL64 0 -6.40890777433692e-21

* Branch 65
Rabr65 node_1 netRa65 5320586.8535108045
Lbr65 netRa65 netL65 -6.128498833526046e-10
Rbbr65 netL65 0 -5557314.28546816
Cbr65 netL65 0 -2.072563112061275e-23

* Branch 66
Rabr66 node_1 netRa66 267175.97810571216
Lbr66 netRa66 netL66 -5.208348958380209e-10
Rbbr66 netL66 0 -2155599.435748113
Cbr66 netL66 0 -9.036019677424607e-22

* Branch 67
Rabr67 node_1 netRa67 947735.1913572169
Lbr67 netRa67 netL67 -7.252488241685864e-10
Rbbr67 netL67 0 -1874893.0413499624
Cbr67 netL67 0 -4.0802205151604613e-22

* Branch 68
Rabr68 node_1 netRa68 2703576.0978250443
Lbr68 netRa68 netL68 7.484999103716268e-10
Rbbr68 netL68 0 -3384872.387863306
Cbr68 netL68 0 8.179894729669515e-23

* Branch 69
Rabr69 node_1 netRa69 5635474.6886766935
Lbr69 netRa69 netL69 -1.8653869893047964e-09
Rbbr69 netL69 0 -6755106.196060356
Cbr69 netL69 0 -4.8996767485501903e-23

* Branch 70
Rabr70 node_1 netRa70 -30388141.007169288
Lbr70 netRa70 netL70 2.610821214806339e-09
Rbbr70 netL70 0 30961383.969140954
Cbr70 netL70 0 2.774874298090518e-24

* Branch 71
Rabr71 node_1 netRa71 3801709.126320424
Lbr71 netRa71 netL71 7.533842018346412e-10
Rbbr71 netL71 0 -4263985.39285041
Cbr71 netL71 0 4.647680292771172e-23

* Branch 72
Rabr72 node_1 netRa72 -3078539.935376403
Lbr72 netRa72 netL72 3.698373662372214e-09
Rbbr72 netL72 0 5146904.102048755
Cbr72 netL72 0 2.3338069346414503e-22

* Branch 73
Rabr73 node_1 netRa73 -1469586.762041098
Lbr73 netRa73 netL73 7.356258935794854e-10
Rbbr73 netL73 0 1885073.1080893
Cbr73 netL73 0 2.655314045102574e-22

* Branch 74
Rabr74 node_1 netRa74 -59877.94150891765
Lbr74 netRa74 netL74 -2.781879826494734e-10
Rbbr74 netL74 0 1557864.9295115522
Cbr74 netL74 0 -2.9831794705260252e-21

* Branch 75
Rabr75 node_1 netRa75 -206244.33745652813
Lbr75 netRa75 netL75 -1.8333829119184884e-10
Rbbr75 netL75 0 334085.08160097187
Cbr75 netL75 0 -2.6609470145097643e-21

* Branch 76
Rabr76 node_1 netRa76 700752.1583067087
Lbr76 netRa76 netL76 -7.226446732323348e-10
Rbbr76 netL76 0 -2162251.267776109
Cbr76 netL76 0 -4.7690173488358115e-22

* Branch 77
Rabr77 node_1 netRa77 150730.3863480556
Lbr77 netRa77 netL77 2.920724526608969e-10
Rbbr77 netL77 0 -1867753.3109711672
Cbr77 netL77 0 1.0375602004685248e-21

* Branch 78
Rabr78 node_1 netRa78 -35735.31948154068
Lbr78 netRa78 netL78 -2.0843709609893267e-10
Rbbr78 netL78 0 1354769.1378413816
Cbr78 netL78 0 -4.306527302582568e-21

* Branch 79
Rabr79 node_1 netRa79 -23541087.388619483
Lbr79 netRa79 netL79 1.998348884217904e-08
Rbbr79 netL79 0 31027913.50136867
Cbr79 netL79 0 2.7358144431764215e-23

* Branch 80
Rabr80 node_1 netRa80 4209437.445119078
Lbr80 netRa80 netL80 1.88048028369076e-08
Rbbr80 netL80 0 -39309390.72825826
Cbr80 netL80 0 1.1365022561949696e-22

* Branch 81
Rabr81 node_1 netRa81 1655640.5893897659
Lbr81 netRa81 netL81 6.1204161021194855e-09
Rbbr81 netL81 0 -10591547.648711266
Cbr81 netL81 0 3.49062200377657e-22

* Branch 82
Rabr82 node_1 netRa82 20482.54830879247
Lbr82 netRa82 netL82 -2.2489614907553218e-10
Rbbr82 netL82 0 -2605350.3120083027
Cbr82 netL82 0 -4.212755058469714e-21

* Branch 83
Rabr83 node_1 netRa83 -15187.151486997152
Lbr83 netRa83 netL83 -4.887754019313526e-11
Rbbr83 netL83 0 208584.91916933536
Cbr83 netL83 0 -1.5431943159719295e-20

* Branch 84
Rabr84 node_1 netRa84 83539.95645640964
Lbr84 netRa84 netL84 -2.165005900455121e-10
Rbbr84 netL84 0 -572427.3359973856
Cbr84 netL84 0 -4.526408893057722e-21

* Branch 85
Rabr85 node_1 netRa85 441.4037018491502
Lbr85 netRa85 netL85 -6.914033024094412e-11
Rbbr85 netL85 0 -14439713.407512099
Cbr85 netL85 0 -1.0711297452910255e-20

* Branch 86
Rabr86 node_1 netRa86 -224806.05658735282
Lbr86 netRa86 netL86 -2.5106338398413245e-10
Rbbr86 netL86 0 878006.122217567
Cbr86 netL86 0 -1.2721131498309605e-21

* Branch 87
Rabr87 node_1 netRa87 -62173.15784497324
Lbr87 netRa87 netL87 -2.0088209674985753e-10
Rbbr87 netL87 0 918371.0572512114
Cbr87 netL87 0 -3.519433990729629e-21

* Branch 88
Rabr88 node_1 netRa88 146128.186480943
Lbr88 netRa88 netL88 -2.665556566846393e-10
Rbbr88 netL88 0 -620095.3377592135
Cbr88 netL88 0 -2.941079754009967e-21

* Branch 89
Rabr89 node_1 netRa89 -9923290.685288822
Lbr89 netRa89 netL89 -1.236102059547763e-09
Rbbr89 netL89 0 10352627.032012861
Cbr89 netL89 0 -1.2032493040211626e-23

* Branch 90
Rabr90 node_1 netRa90 11607565.729199834
Lbr90 netRa90 netL90 -1.0878918438468245e-09
Rbbr90 netL90 0 -11897735.077337265
Cbr90 netL90 0 -7.877247829943124e-24

* Branch 91
Rabr91 node_1 netRa91 78717.60088933689
Lbr91 netRa91 netL91 -2.15176567901104e-10
Rbbr91 netL91 0 -672840.8855576135
Cbr91 netL91 0 -4.061052342812589e-21

* Branch 92
Rabr92 node_1 netRa92 41055.642042061576
Lbr92 netRa92 netL92 -1.4105731471505573e-10
Rbbr92 netL92 0 -359262.0090251191
Cbr92 netL92 0 -9.557135250229236e-21

* Branch 93
Rabr93 node_1 netRa93 40303.62661088609
Lbr93 netRa93 netL93 -1.1429091560650535e-10
Rbbr93 netL93 0 -521371.08161690395
Cbr93 netL93 0 -5.435026122122333e-21

* Branch 94
Rabr94 node_1 netRa94 -21078.93597959106
Lbr94 netRa94 netL94 -1.5225224579127047e-10
Rbbr94 netL94 0 1225261.3760820818
Cbr94 netL94 0 -5.906282162429696e-21

* Branch 95
Rabr95 node_1 netRa95 -3241839.797899396
Lbr95 netRa95 netL95 -7.522139401394645e-10
Rbbr95 netL95 0 3400290.8707892983
Cbr95 netL95 0 -6.824760234506312e-23

* Branch 96
Rabr96 node_1 netRa96 -249035.82942351248
Lbr96 netRa96 netL96 -1.8609520452011853e-10
Rbbr96 netL96 0 366197.95665562846
Cbr96 netL96 0 -2.0415874056229956e-21

* Branch 97
Rabr97 node_1 netRa97 -1286709.1994865923
Lbr97 netRa97 netL97 -4.487162035570832e-10
Rbbr97 netL97 0 1434321.1653349625
Cbr97 netL97 0 -2.431888475983513e-22

* Branch 98
Rabr98 node_1 netRa98 -358234.6736436552
Lbr98 netRa98 netL98 -1.9971070897263342e-10
Rbbr98 netL98 0 448651.83796094527
Cbr98 netL98 0 -1.2431745032028342e-21

* Branch 99
Rabr99 node_1 netRa99 -163361.44895187105
Lbr99 netRa99 netL99 1.6178792294417613e-10
Rbbr99 netL99 0 355922.4704263336
Cbr99 netL99 0 2.7792859655106804e-21

.ends


* Y'12
.subckt yp12 node_1 node_2
* Branch 0
Rabr0 node_1 netRa0 -4548.329385620524
Lbr0 netRa0 netL0 -8.61879320682396e-12
Rbbr0 netL0 node_2 37144.25992410874
Cbr0 netL0 node_2 -1.0269269499876077e-19

* Branch 1
Rabr1 node_1 netRa1 -9655.547703585782
Lbr1 netRa1 netL1 -9.421451827577144e-12
Rbbr1 netL1 node_2 21258.612168012427
Cbr1 netL1 node_2 -6.106968841814993e-20

* Branch 2
Rabr2 node_1 netRa2 -2463.1131037610207
Lbr2 netRa2 netL2 -6.820460619888718e-12
Rbbr2 netL2 node_2 61864.411209089616
Cbr2 netL2 node_2 -1.397112680939911e-19

* Branch 3
Rabr3 node_1 netRa3 -143.79156608009507
Lbr3 netRa3 netL3 -4.81927251240386e-12
Rbbr3 netL3 node_2 -28095.957121885687
Cbr3 netL3 node_2 -1.9640687787542967e-19

* Branch 4
Rabr4 node_1 netRa4 450.4790643502964
Lbr4 netRa4 netL4 -2.7353233037655358e-12
Rbbr4 netL4 node_2 -12364.039594847836
Cbr4 netL4 node_2 -3.089517634664347e-19

* Branch 5
Rabr5 node_1 netRa5 -2068.8762582919026
Lbr5 netRa5 netL5 2.8508711751435124e-12
Rbbr5 netL5 node_2 13604.929480113527
Cbr5 netL5 node_2 9.623091486350787e-20

* Branch 6
Rabr6 node_1 netRa6 -2217.695878284633
Lbr6 netRa6 netL6 1.4046863597812456e-12
Rbbr6 netL6 node_2 4908.971732231919
Cbr6 netL6 node_2 1.265472676248742e-19

* Branch 7
Rabr7 node_1 netRa7 795.1662785060912
Lbr7 netRa7 netL7 1.1648812690625122e-12
Rbbr7 netL7 node_2 -4290.58267023373
Cbr7 netL7 node_2 3.574669882471934e-19

* Branch 8
Rabr8 node_1 netRa8 12051.621848166997
Lbr8 netRa8 netL8 3.952273945531996e-12
Rbbr8 netL8 node_2 -16703.02702866692
Cbr8 netL8 node_2 1.9827380326043002e-20

* Branch 9
Rabr9 node_1 netRa9 -3191.720117214
Lbr9 netRa9 netL9 -1.3681097241587631e-12
Rbbr9 netL9 node_2 5226.351743233781
Cbr9 netL9 node_2 -8.29849256327212e-20

* Branch 10
Rabr10 node_1 netRa10 1238.0297759023852
Lbr10 netRa10 netL10 -1.890631433349891e-12
Rbbr10 netL10 node_2 -4990.023400921194
Cbr10 netL10 node_2 -2.9438215806905185e-19

* Branch 11
Rabr11 node_1 netRa11 442.87743237809826
Lbr11 netRa11 netL11 9.28461593657386e-13
Rbbr11 netL11 node_2 -4467.272987853787
Cbr11 netL11 node_2 4.962502238183596e-19

* Branch 12
Rabr12 node_1 netRa12 -31551.594372565494
Lbr12 netRa12 netL12 3.4583760281750825e-12
Rbbr12 netL12 node_2 32721.074698082262
Cbr12 netL12 node_2 3.3404728431809807e-21

* Branch 13
Rabr13 node_1 netRa13 1169.816611479573
Lbr13 netRa13 netL13 -6.05254712565486e-12
Rbbr13 netL13 node_2 -13153.237669257307
Cbr13 netL13 node_2 -3.513013570776874e-19

* Branch 14
Rabr14 node_1 netRa14 1763.3197571357787
Lbr14 netRa14 netL14 -6.040645552591912e-13
Rbbr14 netL14 node_2 -2407.798713193065
Cbr14 netL14 node_2 -1.4119515523443436e-19

* Branch 15
Rabr15 node_1 netRa15 8809.10034957307
Lbr15 netRa15 netL15 -1.5813296537556295e-12
Rbbr15 netL15 node_2 -9545.548860024473
Cbr15 netL15 node_2 -1.8730989407487576e-20

* Branch 16
Rabr16 node_1 netRa16 6080.620655815042
Lbr16 netRa16 netL16 8.085721095571799e-13
Rbbr16 netL16 node_2 -6398.268523663684
Cbr16 netL16 node_2 2.0838087284737143e-20

* Branch 17
Rabr17 node_1 netRa17 -765.5258771862933
Lbr17 netRa17 netL17 1.0616243991014298e-12
Rbbr17 netL17 node_2 3585.6450806659313
Cbr17 netL17 node_2 3.765658745894417e-19

* Branch 18
Rabr18 node_1 netRa18 3315.6684306415937
Lbr18 netRa18 netL18 -1.3634316189247533e-12
Rbbr18 netL18 node_2 -4659.413394276335
Cbr18 netL18 node_2 -8.762416629764239e-20

* Branch 19
Rabr19 node_1 netRa19 930.4850628267898
Lbr19 netRa19 netL19 6.823857285497428e-13
Rbbr19 netL19 node_2 -2356.775718789886
Cbr19 netL19 node_2 3.1473241307932497e-19

* Branch 20
Rabr20 node_1 netRa20 20104.305544873343
Lbr20 netRa20 netL20 6.918869057153328e-12
Rbbr20 netL20 node_2 -25588.970900860953
Cbr20 netL20 node_2 1.351973435473039e-20

* Branch 21
Rabr21 node_1 netRa21 -2089.1679873645458
Lbr21 netRa21 netL21 -4.412672913292193e-12
Rbbr21 netL21 node_2 6374.314388226705
Cbr21 netL21 node_2 -3.418283387852535e-19

* Branch 22
Rabr22 node_1 netRa22 670.8690582261719
Lbr22 netRa22 netL22 -1.0497371398543144e-12
Rbbr22 netL22 node_2 -5821.211298126784
Cbr22 netL22 node_2 -2.6306824892804503e-19

* Branch 23
Rabr23 node_1 netRa23 184.71108363805214
Lbr23 netRa23 netL23 4.605450878787348e-13
Rbbr23 netL23 node_2 -3633.1091117532865
Cbr23 netL23 node_2 7.109036513308015e-19

* Branch 24
Rabr24 node_1 netRa24 28927.432438034484
Lbr24 netRa24 netL24 -3.485146595619764e-12
Rbbr24 netL24 node_2 -29690.00557509124
Cbr24 netL24 node_2 -4.0516432472923736e-21

* Branch 25
Rabr25 node_1 netRa25 912228.8076180632
Lbr25 netRa25 netL25 1.4454350266363379e-11
Rbbr25 netL25 node_2 -912851.8160170903
Cbr25 netL25 node_2 1.7361106151076064e-23

* Branch 26
Rabr26 node_1 netRa26 3832.6231077181856
Lbr26 netRa26 netL26 -1.8672974369125225e-12
Rbbr26 netL26 node_2 -5344.682056605138
Cbr26 netL26 node_2 -9.070196963316938e-20

* Branch 27
Rabr27 node_1 netRa27 3001.5010737458756
Lbr27 netRa27 netL27 -9.63370702739997e-13
Rbbr27 netL27 node_2 -3945.992879656781
Cbr27 netL27 node_2 -8.10722421722952e-20

* Branch 28
Rabr28 node_1 netRa28 -8361.608640300401
Lbr28 netRa28 netL28 -1.094031360359582e-12
Rbbr28 netL28 node_2 8843.071025981866
Cbr28 netL28 node_2 -1.4815067068953e-20

* Branch 29
Rabr29 node_1 netRa29 2934.938294898914
Lbr29 netRa29 netL29 -1.144049604896681e-12
Rbbr29 netL29 node_2 -3929.089805839541
Cbr29 netL29 node_2 -9.885465959666894e-20

* Branch 30
Rabr30 node_1 netRa30 3024.6510217709097
Lbr30 netRa30 netL30 1.143788560014836e-12
Rbbr30 netL30 node_2 -3897.407224909318
Cbr30 netL30 node_2 9.736424402293913e-20

* Branch 31
Rabr31 node_1 netRa31 -1350.1117856183619
Lbr31 netRa31 netL31 -2.899462666123085e-12
Rbbr31 netL31 node_2 4324.632139789816
Cbr31 netL31 node_2 -5.065120823886234e-19

* Branch 32
Rabr32 node_1 netRa32 2291.600546906324
Lbr32 netRa32 netL32 -8.625082703641023e-13
Rbbr32 netL32 node_2 -3258.9380180711546
Cbr32 netL32 node_2 -1.1510393839336306e-19

* Branch 33
Rabr33 node_1 netRa33 938.3801672085297
Lbr33 netRa33 netL33 -1.7736413494529754e-12
Rbbr33 netL33 node_2 -5232.118874548823
Cbr33 netL33 node_2 -3.555321822834436e-19

* Branch 34
Rabr34 node_1 netRa34 2918.125217014603
Lbr34 netRa34 netL34 -1.4116820186934115e-12
Rbbr34 netL34 node_2 -4404.852632618594
Cbr34 netL34 node_2 -1.093770721130527e-19

* Branch 35
Rabr35 node_1 netRa35 25660.35112128309
Lbr35 netRa35 netL35 6.131606969168549e-12
Rbbr35 netL35 node_2 -30489.01649504496
Cbr35 netL35 node_2 7.853186098092487e-21

* Branch 36
Rabr36 node_1 netRa36 2761.759553351607
Lbr36 netRa36 netL36 -1.9254468706733945e-12
Rbbr36 netL36 node_2 -4802.955366049448
Cbr36 netL36 node_2 -1.4455011737671225e-19

* Branch 37
Rabr37 node_1 netRa37 11545.17471694387
Lbr37 netRa37 netL37 4.004866866978394e-12
Rbbr37 netL37 node_2 -15009.642824538145
Cbr37 netL37 node_2 2.3148778001368643e-20

* Branch 38
Rabr38 node_1 netRa38 29947.978651588288
Lbr38 netRa38 netL38 5.540673006447626e-12
Rbbr38 netL38 node_2 -32062.89592278224
Cbr38 netL38 node_2 5.774431467422203e-21

* Branch 39
Rabr39 node_1 netRa39 -69781.33155756039
Lbr39 netRa39 netL39 -2.4997683414682596e-11
Rbbr39 netL39 node_2 78542.51119948283
Cbr39 netL39 node_2 -4.566666304117486e-21

* Branch 40
Rabr40 node_1 netRa40 1854.9974403264089
Lbr40 netRa40 netL40 -3.5779870355678027e-12
Rbbr40 netL40 node_2 -10062.711989360141
Cbr40 netL40 node_2 -1.905485142159522e-19

* Branch 41
Rabr41 node_1 netRa41 -2270.1818234436496
Lbr41 netRa41 netL41 -2.7756942060061437e-12
Rbbr41 netL41 node_2 3938.296239449046
Cbr41 netL41 node_2 -3.1160773301653963e-19

* Branch 42
Rabr42 node_1 netRa42 -58237233.36473126
Lbr42 netRa42 netL42 4.617573316720905e-10
Rbbr42 netL42 node_2 58239417.79877633
Cbr42 netL42 node_2 1.3614132259948444e-25

* Branch 43
Rabr43 node_1 netRa43 -7945.577809921136
Lbr43 netRa43 netL43 -4.492751789624777e-12
Rbbr43 netL43 node_2 12704.598783039859
Cbr43 netL43 node_2 -4.4547651416290276e-20

* Branch 44
Rabr44 node_1 netRa44 -26194.628130484532
Lbr44 netRa44 netL44 -8.08971445177033e-12
Rbbr44 netL44 node_2 30984.44828038505
Cbr44 netL44 node_2 -9.97179431327881e-21

* Branch 45
Rabr45 node_1 netRa45 -163977869.98222342
Lbr45 netRa45 netL45 -7.482479982630111e-10
Rbbr45 netL45 node_2 163979728.06773147
Cbr45 netL45 node_2 -2.7827398787151336e-26

* Branch 46
Rabr46 node_1 netRa46 -108691.47812288617
Lbr46 netRa46 netL46 1.7567271237138848e-11
Rbbr46 netL46 node_2 110308.74270075573
Cbr46 netL46 node_2 1.4649184968221005e-21

* Branch 47
Rabr47 node_1 netRa47 -7607.037629579046
Lbr47 netRa47 netL47 8.036698425819759e-12
Rbbr47 netL47 node_2 27369.50933265488
Cbr47 netL47 node_2 3.856282521197166e-20

* Branch 48
Rabr48 node_1 netRa48 -1173.5695947717609
Lbr48 netRa48 netL48 -2.0827695037462454e-12
Rbbr48 netL48 node_2 4473.690880970327
Cbr48 netL48 node_2 -3.971499918068684e-19

* Branch 49
Rabr49 node_1 netRa49 11178.182503010901
Lbr49 netRa49 netL49 -4.8784152915927695e-12
Rbbr49 netL49 node_2 -15673.91591330491
Cbr49 netL49 node_2 -2.78373830572262e-20

* Branch 50
Rabr50 node_1 netRa50 102161.39414998714
Lbr50 netRa50 netL50 1.9705700626506336e-11
Rbbr50 netL50 node_2 -111861.88372053792
Cbr50 netL50 node_2 1.7245168928374325e-21

* Branch 51
Rabr51 node_1 netRa51 -322906.6352398361
Lbr51 netRa51 netL51 -3.491031465317884e-11
Rbbr51 netL51 node_2 325373.3144189109
Cbr51 netL51 node_2 -3.322892792082444e-22

* Branch 52
Rabr52 node_1 netRa52 -67253.93976588252
Lbr52 netRa52 netL52 -1.4871079570366144e-11
Rbbr52 netL52 node_2 69500.45660907478
Cbr52 netL52 node_2 -3.1818504648161447e-21

* Branch 53
Rabr53 node_1 netRa53 -28255.971167706448
Lbr53 netRa53 netL53 5.147033617839698e-12
Rbbr53 netL53 node_2 28774.38324651601
Cbr53 netL53 node_2 6.330103410661101e-21

* Branch 54
Rabr54 node_1 netRa54 -166705.7408039627
Lbr54 netRa54 netL54 -1.9543208880378082e-11
Rbbr54 netL54 node_2 168137.22980327928
Cbr54 netL54 node_2 -6.972668484444149e-22

* Branch 55
Rabr55 node_1 netRa55 -28906.826387615463
Lbr55 netRa55 netL55 -5.252673856734171e-12
Rbbr55 netL55 node_2 29499.689257934577
Cbr55 netL55 node_2 -6.160085365636105e-21

* Branch 56
Rabr56 node_1 netRa56 -8445.388279767842
Lbr56 netRa56 netL56 -4.91536400659729e-12
Rbbr56 netL56 node_2 10574.376986246134
Cbr56 netL56 node_2 -5.50412716810764e-20

* Branch 57
Rabr57 node_1 netRa57 -12229.5386864159
Lbr57 netRa57 netL57 -6.380000607318893e-12
Rbbr57 netL57 node_2 14811.276618150045
Cbr57 netL57 node_2 -3.522293648160867e-20

* Branch 58
Rabr58 node_1 netRa58 -105713.27656430738
Lbr58 netRa58 netL58 -1.9850876102440796e-11
Rbbr58 netL58 node_2 108371.98892452293
Cbr58 netL58 node_2 -1.7327552072936467e-21

* Branch 59
Rabr59 node_1 netRa59 42118.315229026266
Lbr59 netRa59 netL59 1.4768597169546983e-11
Rbbr59 netL59 node_2 -55633.58258713719
Cbr59 netL59 node_2 6.303047730698847e-21

* Branch 60
Rabr60 node_1 netRa60 -56601.2413592831
Lbr60 netRa60 netL60 -1.3374600431137199e-11
Rbbr60 netL60 node_2 59256.9417017971
Cbr60 netL60 node_2 -3.987853409161506e-21

* Branch 61
Rabr61 node_1 netRa61 -3942.642681552307
Lbr61 netRa61 netL61 -2.4542575277778537e-12
Rbbr61 netL61 node_2 5064.222481636241
Cbr61 netL61 node_2 -1.2293696835320373e-19

* Branch 62
Rabr62 node_1 netRa62 55399.0152253681
Lbr62 netRa62 netL62 -1.0990113559714508e-11
Rbbr62 netL62 node_2 -60589.79059865117
Cbr62 netL62 node_2 -3.2740041998989787e-21

* Branch 63
Rabr63 node_1 netRa63 -8221.096001701464
Lbr63 netRa63 netL63 -4.647716498624117e-12
Rbbr63 netL63 node_2 10697.648008977805
Cbr63 netL63 node_2 -5.285475936101531e-20

* Branch 64
Rabr64 node_1 netRa64 -100191.81402443028
Lbr64 netRa64 netL64 -1.7697976119029496e-11
Rbbr64 netL64 node_2 102716.58548475387
Cbr64 netL64 node_2 -1.7197709681664273e-21

* Branch 65
Rabr65 node_1 netRa65 -9522.586202758184
Lbr65 netRa65 netL65 4.281258066575199e-12
Rbbr65 netL65 node_2 10522.363733235283
Cbr65 netL65 node_2 4.272095274385937e-20

* Branch 66
Rabr66 node_1 netRa66 -6896.840535493026
Lbr66 netRa66 netL66 -3.97467546908344e-12
Rbbr66 netL66 node_2 8977.82770293403
Cbr66 netL66 node_2 -6.420462334870424e-20

* Branch 67
Rabr67 node_1 netRa67 29865.47026363689
Lbr67 netRa67 netL67 1.1118167916056999e-11
Rbbr67 netL67 node_2 -40909.272087038225
Cbr67 netL67 node_2 9.101198724966172e-21

* Branch 68
Rabr68 node_1 netRa68 5486.825527804837
Lbr68 netRa68 netL68 2.1683099916878998e-11
Rbbr68 netL68 node_2 -129703.63939219169
Cbr68 netL68 node_2 3.051763062661189e-20

* Branch 69
Rabr69 node_1 netRa69 160244.62868527343
Lbr69 netRa69 netL69 2.2607239891240325e-11
Rbbr69 netL69 node_2 -168018.76265958822
Cbr69 netL69 node_2 8.39716593464522e-22

* Branch 70
Rabr70 node_1 netRa70 -585.2201493289308
Lbr70 netRa70 netL70 2.2550616647961666e-12
Rbbr70 netL70 node_2 24218.22551438981
Cbr70 netL70 node_2 1.5883210081570768e-19

* Branch 71
Rabr71 node_1 netRa71 111363.25682352175
Lbr71 netRa71 netL71 2.2638281724136173e-11
Rbbr71 netL71 node_2 -119479.22196886614
Cbr71 netL71 node_2 1.7015965162739206e-21

* Branch 72
Rabr72 node_1 netRa72 1141.0080088125374
Lbr72 netRa72 netL72 1.358212194771603e-11
Rbbr72 netL72 node_2 -265611.6225590392
Cbr72 netL72 node_2 4.5105389081528786e-20

* Branch 73
Rabr73 node_1 netRa73 9369.772171677727
Lbr73 netRa73 netL73 1.3794652260839063e-11
Rbbr73 netL73 node_2 -39669.77818594612
Cbr73 netL73 node_2 3.714451485368332e-20

* Branch 74
Rabr74 node_1 netRa74 -153542.79579982092
Lbr74 netRa74 netL74 2.7548118249661995e-11
Rbbr74 netL74 node_2 162508.6701433469
Cbr74 netL74 node_2 1.1039264022553096e-21

* Branch 75
Rabr75 node_1 netRa75 -15333.182284208991
Lbr75 netRa75 netL75 7.473641964303426e-12
Rbbr75 netL75 node_2 18514.020987032014
Cbr75 netL75 node_2 2.6318920902801983e-20

* Branch 76
Rabr76 node_1 netRa76 17470.937270729522
Lbr76 netRa76 netL76 1.4390795632009187e-11
Rbbr76 netL76 node_2 -37839.61427148141
Cbr76 netL76 node_2 2.1780066546693356e-20

* Branch 77
Rabr77 node_1 netRa77 -5125.553881341777
Lbr77 netRa77 netL77 5.0847316691456426e-12
Rbbr77 netL77 node_2 10225.061736044674
Cbr77 netL77 node_2 9.695225351508071e-20

* Branch 78
Rabr78 node_1 netRa78 -5342.305207799958
Lbr78 netRa78 netL78 5.22448772802774e-12
Rbbr78 netL78 node_2 10693.762862791938
Cbr78 netL78 node_2 9.138651452738664e-20

* Branch 79
Rabr79 node_1 netRa79 29764.679933934123
Lbr79 netRa79 netL79 1.733774630185483e-11
Rbbr79 netL79 node_2 -45718.72691793301
Cbr79 netL79 node_2 1.2746286600659747e-20

* Branch 80
Rabr80 node_1 netRa80 10825.120334926005
Lbr80 netRa80 netL80 1.0300428175054345e-11
Rbbr80 netL80 node_2 -23373.331284794273
Cbr80 netL80 node_2 4.073904467399371e-20

* Branch 81
Rabr81 node_1 netRa81 365729.48340259294
Lbr81 netRa81 netL81 2.496281507114599e-11
Rbbr81 netL81 node_2 -369419.7130049154
Cbr81 netL81 node_2 1.8477196350238562e-22

* Branch 82
Rabr82 node_1 netRa82 -8731.704572312334
Lbr82 netRa82 netL82 5.869564752235954e-12
Rbbr82 netL82 node_2 13012.445217061379
Cbr82 netL82 node_2 5.163223198063753e-20

* Branch 83
Rabr83 node_1 netRa83 6381.624894643002
Lbr83 netRa83 netL83 7.619572426169391e-12
Rbbr83 netL83 node_2 -16950.0196301232
Cbr83 netL83 node_2 7.051640886426414e-20

* Branch 84
Rabr84 node_1 netRa84 2796.7583114329905
Lbr84 netRa84 netL84 6.260685116296532e-12
Rbbr84 netL84 node_2 -20200.462724091343
Cbr84 netL84 node_2 1.1104456812335005e-19

* Branch 85
Rabr85 node_1 netRa85 -10848.32454416493
Lbr85 netRa85 netL85 -3.651731883333941e-12
Rbbr85 netL85 node_2 11670.040136359923
Cbr85 netL85 node_2 -2.885350640939421e-20

* Branch 86
Rabr86 node_1 netRa86 2231.7480493523385
Lbr86 netRa86 netL86 5.339058077448903e-12
Rbbr86 netL86 node_2 -16598.182664594842
Cbr86 netL86 node_2 1.444558909919985e-19

* Branch 87
Rabr87 node_1 netRa87 10091.45534091619
Lbr87 netRa87 netL87 8.517691836322298e-12
Rbbr87 netL87 node_2 -20191.89936813531
Cbr87 netL87 node_2 4.1835527066712897e-20

* Branch 88
Rabr88 node_1 netRa88 3799.4990334378085
Lbr88 netRa88 netL88 6.164335424027626e-12
Rbbr88 netL88 node_2 -17440.775780994485
Cbr88 netL88 node_2 9.317423053981227e-20

* Branch 89
Rabr89 node_1 netRa89 1181.9948646219216
Lbr89 netRa89 netL89 5.036608773802011e-12
Rbbr89 netL89 node_2 -29643.479975509865
Cbr89 netL89 node_2 1.443669855393669e-19

* Branch 90
Rabr90 node_1 netRa90 -3263.6694081543515
Lbr90 netRa90 netL90 5.406565534431014e-12
Rbbr90 netL90 node_2 18208.317533710775
Cbr90 netL90 node_2 9.082303202933253e-20

* Branch 91
Rabr91 node_1 netRa91 -410.99610701853044
Lbr91 netRa91 netL91 5.926457952502622e-12
Rbbr91 netL91 node_2 129418.6410991622
Cbr91 netL91 node_2 1.096091600283929e-19

* Branch 92
Rabr92 node_1 netRa92 5925.255820994423
Lbr92 netRa92 netL92 5.87655145471596e-12
Rbbr92 netL92 node_2 -12918.040234305134
Cbr92 netL92 node_2 7.686782961197611e-20

* Branch 93
Rabr93 node_1 netRa93 -5089.803918308199
Lbr93 netRa93 netL93 3.4388405866099943e-12
Rbbr93 netL93 node_2 7357.866791100724
Cbr93 netL93 node_2 9.174645663573458e-20

* Branch 94
Rabr94 node_1 netRa94 12493.271973254767
Lbr94 netRa94 netL94 3.0605467847016275e-12
Rbbr94 netL94 node_2 -14155.128811331182
Cbr94 netL94 node_2 1.7315965243465246e-20

* Branch 95
Rabr95 node_1 netRa95 -841.4744415344022
Lbr95 netRa95 netL95 1.4135828918161044e-12
Rbbr95 netL95 node_2 7407.598949115433
Cbr95 netL95 node_2 2.252754336597724e-19

* Branch 96
Rabr96 node_1 netRa96 -512.2245202841556
Lbr96 netRa96 netL96 6.047315263438153e-13
Rbbr96 netL96 node_2 866.5122914591159
Cbr96 netL96 node_2 1.3552458812322088e-18

* Branch 97
Rabr97 node_1 netRa97 -254.82219346457637
Lbr97 netRa97 netL97 5.318327904386024e-13
Rbbr97 netL97 node_2 2365.7052282965346
Cbr97 netL97 node_2 8.554278525162161e-19

* Branch 98
Rabr98 node_1 netRa98 4045.598076592841
Lbr98 netRa98 netL98 -6.015649603140623e-13
Rbbr98 netL98 node_2 -4344.333986587868
Cbr98 netL98 node_2 -3.41414561649621e-20

* Branch 99
Rabr99 node_1 netRa99 8060.3405765604975
Lbr99 netRa99 netL99 -3.079360274189755e-12
Rbbr99 netL99 node_2 -11669.75050007407
Cbr99 netL99 node_2 -3.221820130795115e-20

.ends


* Y'22
.subckt yp22 node_2 0
* Branch 0
Rabr0 node_2 netRa0 -26126.304283674202
Lbr0 netRa0 netL0 1.6423055384113456e-11
Rbbr0 netL0 0 48548.309914855665
Cbr0 netL0 0 1.2488696478633102e-20

* Branch 1
Rabr1 node_2 netRa1 -61319.02657588663
Lbr1 netRa1 netL1 2.5433045081087287e-11
Rbbr1 netL1 0 84585.196295483
Cbr1 netL1 0 4.793682023654537e-21

* Branch 2
Rabr2 node_2 netRa2 -464450.7734731441
Lbr2 netRa2 netL2 -7.614934484563921e-11
Rbbr2 netL2 0 492929.78290505224
Cbr2 netL2 0 -3.352862616046092e-22

* Branch 3
Rabr3 node_2 netRa3 -2954508.1709165704
Lbr3 netRa3 netL3 -2.031222034135034e-10
Rbbr3 netL3 0 2974126.9139571567
Cbr3 netL3 0 -2.3191999032738502e-23

* Branch 4
Rabr4 node_2 netRa4 30474.786801210466
Lbr4 netRa4 netL4 3.251963957291942e-11
Rbbr4 netL4 0 -92743.51489675147
Cbr4 netL4 0 1.2116456785444627e-20

* Branch 5
Rabr5 node_2 netRa5 -867571.7665996011
Lbr5 netRa5 netL5 1.139745306277173e-10
Rbbr5 netL5 0 888294.552299478
Cbr5 netL5 0 1.4700477783480045e-22

* Branch 6
Rabr6 node_2 netRa6 -64476.93096062781
Lbr6 netRa6 netL6 -2.669859448346379e-11
Rbbr6 netL6 0 89975.62296812708
Cbr6 netL6 0 -4.691060397729504e-21

* Branch 7
Rabr7 node_2 netRa7 -770840.388707006
Lbr7 netRa7 netL7 9.464061207284951e-11
Rbbr7 netL7 0 786644.9455985235
Cbr7 netL7 0 1.5530220752469013e-22

* Branch 8
Rabr8 node_2 netRa8 19151.693946551386
Lbr8 netRa8 netL8 3.180202411406339e-11
Rbbr8 netL8 0 -115064.6068440164
Cbr8 netL8 0 1.546652910471642e-20

* Branch 9
Rabr9 node_2 netRa9 7855.0056308116
Lbr9 netRa9 netL9 -1.1019492499822391e-11
Rbbr9 netL9 0 -41151.90672057621
Cbr9 netL9 0 -3.226867011936146e-20

* Branch 10
Rabr10 node_2 netRa10 34670.97271155243
Lbr10 netRa10 netL10 3.800828103264128e-11
Rbbr10 netL10 0 -108930.36686852043
Cbr10 netL10 0 1.0519438061100218e-20

* Branch 11
Rabr11 node_2 netRa11 -160648.7504378326
Lbr11 netRa11 netL11 4.6119851991433075e-11
Rbbr11 netL11 0 178896.4857934413
Cbr11 netL11 0 1.5869010863297857e-21

* Branch 12
Rabr12 node_2 netRa12 -94760.67691791347
Lbr12 netRa12 netL12 3.385872070974709e-11
Rbbr12 netL12 0 111419.01366988981
Cbr12 netL12 0 3.164902246686087e-21

* Branch 13
Rabr13 node_2 netRa13 25758.494681690707
Lbr13 netRa13 netL13 4.175292486921247e-11
Rbbr13 netL13 0 -147038.28362607784
Cbr13 netL13 0 1.1628456864086572e-20

* Branch 14
Rabr14 node_2 netRa14 4065.962025941412
Lbr14 netRa14 netL14 3.491048288163835e-12
Rbbr14 netL14 0 -11148.075338843395
Cbr14 netL14 0 7.864117257739037e-20

* Branch 15
Rabr15 node_2 netRa15 85822.82361390526
Lbr15 netRa15 netL15 6.862572309771516e-11
Rbbr15 netL15 0 -182015.11257766304
Cbr15 netL15 0 4.479116832429558e-21

* Branch 16
Rabr16 node_2 netRa16 10814.14415978469
Lbr16 netRa16 netL16 -8.738330132078946e-12
Rbbr16 netL16 0 -20398.880768784285
Cbr16 netL16 0 -3.897507451111352e-20

* Branch 17
Rabr17 node_2 netRa17 212.58152654483985
Lbr17 netRa17 netL17 9.36137391365165e-12
Rbbr17 netL17 0 -5318010.597384953
Cbr17 netL17 0 3.2831990818875885e-20

* Branch 18
Rabr18 node_2 netRa18 95005.70166533632
Lbr18 netRa18 netL18 -4.3536347291267384e-11
Rbbr18 netL18 0 -138523.24395510968
Cbr18 netL18 0 -3.2847786737741196e-21

* Branch 19
Rabr19 node_2 netRa19 16241.145678375493
Lbr19 netRa19 netL19 2.4731075315828416e-11
Rbbr19 netL19 0 -72611.40263404313
Cbr19 netL19 0 2.1412554308614424e-20

* Branch 20
Rabr20 node_2 netRa20 11774.995148567208
Lbr20 netRa20 netL20 -1.2940977494502987e-11
Rbbr20 netL20 0 -47729.997460911356
Cbr20 netL20 0 -2.2691821532890117e-20

* Branch 21
Rabr21 node_2 netRa21 2058.3661118524165
Lbr21 netRa21 netL21 1.4665329025972115e-11
Rbbr21 netL21 0 -83985.3872337311
Cbr21 netL21 0 9.350817852713877e-20

* Branch 22
Rabr22 node_2 netRa22 6641064.421957778
Lbr22 netRa22 netL22 -1.3456607629263527e-10
Rbbr22 netL22 0 -6646514.933657939
Cbr22 netL22 0 -3.047833103525288e-24

* Branch 23
Rabr23 node_2 netRa23 254802.9005794528
Lbr23 netRa23 netL23 -5.806984847266747e-11
Rbbr23 netL23 0 -282186.2536567472
Cbr23 netL23 0 -8.053122219930365e-22

* Branch 24
Rabr24 node_2 netRa24 21489540.74790357
Lbr24 netRa24 netL24 -5.938102361103511e-10
Rbbr24 netL24 0 -21499105.11473774
Cbr24 netL24 0 -1.2848477152110846e-24

* Branch 25
Rabr25 node_2 netRa25 -17431.717342831464
Lbr25 netRa25 netL25 1.3606989038638087e-11
Rbbr25 netL25 0 35002.26552876175
Cbr25 netL25 0 2.2090470738188224e-20

* Branch 26
Rabr26 node_2 netRa26 429417.2172558133
Lbr26 netRa26 netL26 8.687981656142709e-11
Rbbr26 netL26 0 -490779.81926156423
Cbr26 netL26 0 4.1325875248869746e-22

* Branch 27
Rabr27 node_2 netRa27 229359.2116149157
Lbr27 netRa27 netL27 -7.302532055428391e-11
Rbbr27 netL27 0 -278748.8914890023
Cbr27 netL27 0 -1.138055252725096e-21

* Branch 28
Rabr28 node_2 netRa28 33854.55837208988
Lbr28 netRa28 netL28 2.3140661955452018e-11
Rbbr28 netL28 0 -45581.85873005601
Cbr28 netL28 0 1.5108923989006498e-20

* Branch 29
Rabr29 node_2 netRa29 13348.953628397854
Lbr29 netRa29 netL29 1.0477533143364336e-11
Rbbr29 netL29 0 -37497.315845172445
Cbr29 netL29 0 2.1113007090220523e-20

* Branch 30
Rabr30 node_2 netRa30 29379.105239982877
Lbr30 netRa30 netL30 -2.609271375605331e-11
Rbbr30 netL30 0 -46762.27331147666
Cbr30 netL30 0 -1.8811123791928152e-20

* Branch 31
Rabr31 node_2 netRa31 -94856.51364689837
Lbr31 netRa31 netL31 7.901357401115763e-11
Rbbr31 netL31 0 139503.24026371998
Cbr31 netL31 0 5.917717731736737e-21

* Branch 32
Rabr32 node_2 netRa32 4129.824722329985
Lbr32 netRa32 netL32 -8.719766446293177e-12
Rbbr32 netL32 0 -46877.18156575093
Cbr32 netL32 0 -4.4041645359443876e-20

* Branch 33
Rabr33 node_2 netRa33 14047.686093788074
Lbr33 netRa33 netL33 1.3708409116635836e-11
Rbbr33 netL33 0 -38145.12520835137
Cbr33 netL33 0 2.584547728223646e-20

* Branch 34
Rabr34 node_2 netRa34 148446.92001850955
Lbr34 netRa34 netL34 -3.199331161443742e-11
Rbbr34 netL34 0 -171705.14976878391
Cbr34 netL34 0 -1.252530490581254e-21

* Branch 35
Rabr35 node_2 netRa35 -22195.501402649938
Lbr35 netRa35 netL35 3.3362316093675523e-11
Rbbr35 netL35 0 102208.85418369978
Cbr35 netL35 0 1.4493162841648885e-20

* Branch 36
Rabr36 node_2 netRa36 3544.534962294288
Lbr36 netRa36 netL36 1.3518699269015335e-11
Rbbr36 netL36 0 -33718.089877956394
Cbr36 netL36 0 1.172889571345702e-19

* Branch 37
Rabr37 node_2 netRa37 2736.04771036185
Lbr37 netRa37 netL37 -2.0480709475999192e-11
Rbbr37 netL37 0 -362345.4547430624
Cbr37 netL37 0 -1.9466971266927664e-20

* Branch 38
Rabr38 node_2 netRa38 4339.3721134567095
Lbr38 netRa38 netL38 -3.036692213051263e-11
Rbbr38 netL38 0 -648313.2845570779
Cbr38 netL38 0 -1.0215716868378313e-20

* Branch 39
Rabr39 node_2 netRa39 -96896.5787165355
Lbr39 netRa39 netL39 3.315033865494889e-11
Rbbr39 netL39 0 126941.16295773475
Cbr39 netL39 0 2.6877125862977026e-21

* Branch 40
Rabr40 node_2 netRa40 -7152.145323464678
Lbr40 netRa40 netL40 2.428299020377707e-11
Rbbr40 netL40 0 50670.6801873417
Cbr40 netL40 0 6.529324302394124e-20

* Branch 41
Rabr41 node_2 netRa41 -14613.914899403842
Lbr41 netRa41 netL41 1.000179129681696e-11
Rbbr41 netL41 0 33204.76872682391
Cbr41 netL41 0 2.0508566203861875e-20

* Branch 42
Rabr42 node_2 netRa42 -44881.115878219796
Lbr42 netRa42 netL42 2.1045016341869356e-11
Rbbr42 netL42 0 75235.83227531999
Cbr42 netL42 0 6.2114645335903085e-21

* Branch 43
Rabr43 node_2 netRa43 31738.915069046066
Lbr43 netRa43 netL43 2.1153654034407568e-11
Rbbr43 netL43 0 -40850.72309677579
Cbr43 netL43 0 1.6393925380283276e-20

* Branch 44
Rabr44 node_2 netRa44 -49080.96134656257
Lbr44 netRa44 netL44 5.137384275528404e-11
Rbbr44 netL44 0 130990.29513839571
Cbr44 netL44 0 7.933454038079839e-21

* Branch 45
Rabr45 node_2 netRa45 10062458.34420978
Lbr45 netRa45 netL45 -2.991349152264094e-10
Rbbr45 netL45 0 -10070282.611784665
Cbr45 netL45 0 -2.9514296565997106e-24

* Branch 46
Rabr46 node_2 netRa46 -213372832.71681693
Lbr46 netRa46 netL46 -2.6711027200971546e-09
Rbbr46 netL46 0 213399056.4670026
Cbr46 netL46 0 -5.866700842720106e-26

* Branch 47
Rabr47 node_2 netRa47 97343.99550867428
Lbr47 netRa47 netL47 -4.650016846601834e-11
Rbbr47 netL47 0 -125899.45302234337
Cbr47 netL47 0 -3.782659593296933e-21

* Branch 48
Rabr48 node_2 netRa48 171580.19038268275
Lbr48 netRa48 netL48 -8.118088220722053e-11
Rbbr48 netL48 0 -196844.51410910045
Cbr48 netL48 0 -2.396408388827248e-21

* Branch 49
Rabr49 node_2 netRa49 -189764.3141126425
Lbr49 netRa49 netL49 4.822021277751388e-11
Rbbr49 netL49 0 221607.98386468642
Cbr49 netL49 0 1.1448463394112644e-21

* Branch 50
Rabr50 node_2 netRa50 16107.04118595093
Lbr50 netRa50 netL50 -2.3174366012231865e-11
Rbbr50 netL50 0 -46564.125461744356
Cbr50 netL50 0 -3.063490279765055e-20

* Branch 51
Rabr51 node_2 netRa51 -16547.280930018445
Lbr51 netRa51 netL51 2.9199676285567654e-11
Rbbr51 netL51 0 48415.2166651383
Cbr51 netL51 0 3.607026241589023e-20

* Branch 52
Rabr52 node_2 netRa52 35482.9399080595
Lbr52 netRa52 netL52 2.580531475659839e-11
Rbbr52 netL52 0 -44651.54638337525
Cbr52 netL52 0 1.635573458890927e-20

* Branch 53
Rabr53 node_2 netRa53 30988.542054241272
Lbr53 netRa53 netL53 -2.5254423650509627e-11
Rbbr53 netL53 0 -58362.07921864876
Cbr53 netL53 0 -1.3901548492937675e-20

* Branch 54
Rabr54 node_2 netRa54 305528.26732253423
Lbr54 netRa54 netL54 -5.503826281165359e-11
Rbbr54 netL54 0 -313744.5528377424
Cbr54 netL54 0 -5.736145884656793e-22

* Branch 55
Rabr55 node_2 netRa55 131477.64533726452
Lbr55 netRa55 netL55 4.9762115114801215e-11
Rbbr55 netL55 0 -187638.41652641087
Cbr55 netL55 0 2.0210482924005664e-21

* Branch 56
Rabr56 node_2 netRa56 -3768.9704414492826
Lbr56 netRa56 netL56 2.1428891485596624e-11
Rbbr56 netL56 0 99748.19789843982
Cbr56 netL56 0 5.556677976538721e-20

* Branch 57
Rabr57 node_2 netRa57 -7414.26577546588
Lbr57 netRa57 netL57 7.465363579689853e-11
Rbbr57 netL57 0 1140861.8148040308
Cbr57 netL57 0 8.44551843078668e-21

* Branch 58
Rabr58 node_2 netRa58 472569.1887269807
Lbr58 netRa58 netL58 -7.564669915277246e-11
Rbbr58 netL58 0 -487191.87582910125
Cbr58 netL58 0 -3.283355338954831e-22

* Branch 59
Rabr59 node_2 netRa59 -70981.59309413013
Lbr59 netRa59 netL59 1.946760339616073e-11
Rbbr59 netL59 0 86317.88990631986
Cbr59 netL59 0 3.173525338323186e-21

* Branch 60
Rabr60 node_2 netRa60 -13026.757220014519
Lbr60 netRa60 netL60 -3.11356400395603e-11
Rbbr60 netL60 0 195686.76423464873
Cbr60 netL60 0 -1.2340459388107553e-20

* Branch 61
Rabr61 node_2 netRa61 -103918.2196359429
Lbr61 netRa61 netL61 1.0276989498883337e-10
Rbbr61 netL61 0 156251.97146806648
Cbr61 netL61 0 6.302553309972899e-21

* Branch 62
Rabr62 node_2 netRa62 721451.6439398082
Lbr62 netRa62 netL62 1.247452163782222e-10
Rbbr62 netL62 0 -762538.4239802832
Cbr62 netL62 0 2.2691111251942273e-22

* Branch 63
Rabr63 node_2 netRa63 364.61656624492
Lbr63 netRa63 netL63 7.97204485251518e-11
Rbbr63 netL63 0 -103885935.77912302
Cbr63 netL63 0 6.907773408769758e-21

* Branch 64
Rabr64 node_2 netRa64 14383005.933207616
Lbr64 netRa64 netL64 -3.380778328953431e-10
Rbbr64 netL64 0 -14392061.836911099
Cbr64 netL64 0 -1.6331327864898008e-24

* Branch 65
Rabr65 node_2 netRa65 -35854.89423424669
Lbr65 netRa65 netL65 -5.795649286014584e-11
Rbbr65 netL65 0 92433.75300534016
Cbr65 netL65 0 -1.7548531426643486e-20

* Branch 66
Rabr66 node_2 netRa66 15775.527662449158
Lbr66 netRa66 netL66 -2.7076656330968302e-11
Rbbr66 netL66 0 -55196.56124497653
Cbr66 netL66 0 -3.098544296379445e-20

* Branch 67
Rabr67 node_2 netRa67 280631.9632231567
Lbr67 netRa67 netL67 3.5774872238944585e-11
Rbbr67 netL67 0 -285624.34345724713
Cbr67 netL67 0 4.464051849393234e-22

* Branch 68
Rabr68 node_2 netRa68 116846288.78440252
Lbr68 netRa68 netL68 2.5318576559648623e-09
Rbbr68 netL68 0 -116948322.05451003
Cbr68 netL68 0 1.852857803438955e-25

* Branch 69
Rabr69 node_2 netRa69 -31701.855482336116
Lbr69 netRa69 netL69 -1.197331880197723e-10
Rbbr69 netL69 0 254487.24858011637
Cbr69 netL69 0 -1.489929375057196e-20

* Branch 70
Rabr70 node_2 netRa70 235482.29343504237
Lbr70 netRa70 netL70 -7.990932406439044e-11
Rbbr70 netL70 0 -269306.39624078706
Cbr70 netL70 0 -1.259722023436667e-21

* Branch 71
Rabr71 node_2 netRa71 26684.41196788366
Lbr71 netRa71 netL71 -3.2244098452943634e-11
Rbbr71 netL71 0 -117306.72273850416
Cbr71 netL71 0 -1.0291024731998236e-20

* Branch 72
Rabr72 node_2 netRa72 -611177.1580222612
Lbr72 netRa72 netL72 1.9437934308763916e-10
Rbbr72 netL72 0 798631.3200299902
Cbr72 netL72 0 3.98179983445154e-22

* Branch 73
Rabr73 node_2 netRa73 -52007.63263170913
Lbr73 netRa73 netL73 -7.211567574082023e-11
Rbbr73 netL73 0 149640.8966235589
Cbr73 netL73 0 -9.268874286622075e-21

* Branch 74
Rabr74 node_2 netRa74 1260379.6286281454
Lbr74 netRa74 netL74 -1.3077513018423582e-10
Rbbr74 netL74 0 -1276271.1884458757
Cbr74 netL74 0 -8.129657841950157e-23

* Branch 75
Rabr75 node_2 netRa75 -128660.02819201114
Lbr75 netRa75 netL75 -3.311754049920183e-10
Rbbr75 netL75 0 2769171.8656140394
Cbr75 netL75 0 -9.298180970467192e-22

* Branch 76
Rabr76 node_2 netRa76 -138866.9848885865
Lbr76 netRa76 netL76 1.8427989314714675e-09
Rbbr76 netL76 0 11513186.746214861
Cbr76 netL76 0 1.1516657636540265e-21

* Branch 77
Rabr77 node_2 netRa77 146873.23330585286
Lbr77 netRa77 netL77 -1.5629553826802977e-10
Rbbr77 netL77 0 -327192.4144869637
Cbr77 netL77 0 -3.2522958580063647e-21

* Branch 78
Rabr78 node_2 netRa78 3311891.918611407
Lbr78 netRa78 netL78 1.4755817427900007e-09
Rbbr78 netL78 0 -3601908.587222307
Cbr78 netL78 0 1.2369615619384895e-22

* Branch 79
Rabr79 node_2 netRa79 4049303.545798885
Lbr79 netRa79 netL79 1.306486519525765e-09
Rbbr79 netL79 0 -4225296.518196758
Cbr79 netL79 0 7.636060578021242e-23

* Branch 80
Rabr80 node_2 netRa80 -164578.82572281544
Lbr80 netRa80 netL80 -2.7612659473932627e-10
Rbbr80 netL80 0 1073364.832356915
Cbr80 netL80 0 -1.5631462471029514e-21

* Branch 81
Rabr81 node_2 netRa81 4401811.005400456
Lbr81 netRa81 netL81 1.2828641047480503e-09
Rbbr81 netL81 0 -4549347.772218734
Cbr81 netL81 0 6.406257475045948e-23

* Branch 82
Rabr82 node_2 netRa82 598185.5899454976
Lbr82 netRa82 netL82 -6.633139926114335e-11
Rbbr82 netL82 0 -605989.1716832939
Cbr82 netL82 0 -1.8298549670375284e-22

* Branch 83
Rabr83 node_2 netRa83 -87919.21235308582
Lbr83 netRa83 netL83 -1.7777433315908985e-10
Rbbr83 netL83 0 401372.2466523917
Cbr83 netL83 0 -5.0382553513278754e-21

* Branch 84
Rabr84 node_2 netRa84 70688.61736347491
Lbr84 netRa84 netL84 -3.0382955049047056e-11
Rbbr84 netL84 0 -83675.6823788027
Cbr84 netL84 0 -5.136518844881521e-21

* Branch 85
Rabr85 node_2 netRa85 -13549.400226577653
Lbr85 netRa85 netL85 1.712538663368889e-11
Rbbr85 netL85 0 56934.181203534354
Cbr85 netL85 0 2.219479263596762e-20

* Branch 86
Rabr86 node_2 netRa86 -336375.1752997769
Lbr86 netRa86 netL86 -1.6834334120580418e-10
Rbbr86 netL86 0 424665.6412308696
Cbr86 netL86 0 -1.1786071998083154e-21

* Branch 87
Rabr87 node_2 netRa87 -10139.507952103411
Lbr87 netRa87 netL87 9.273174197046737e-12
Rbbr87 netL87 0 33565.60029407082
Cbr87 netL87 0 2.7240057980954365e-20

* Branch 88
Rabr88 node_2 netRa88 -10264.280639919456
Lbr88 netRa88 netL88 -3.1387431753177194e-11
Rbbr88 netL88 0 325631.05317016516
Cbr88 netL88 0 -9.40041430420393e-21

* Branch 89
Rabr89 node_2 netRa89 395149.0250143957
Lbr89 netRa89 netL89 -1.2721721075520435e-10
Rbbr89 netL89 0 -509318.9370664543
Cbr89 netL89 0 -6.320368285473903e-22

* Branch 90
Rabr90 node_2 netRa90 -16562.683633434208
Lbr90 netRa90 netL90 -2.384315950450811e-11
Rbbr90 netL90 0 49420.806337709866
Cbr90 netL90 0 -2.914502141814838e-20

* Branch 91
Rabr91 node_2 netRa91 -82539.9081162245
Lbr91 netRa91 netL91 -6.821974895761096e-11
Rbbr91 netL91 0 271828.19816356525
Cbr91 netL91 0 -3.041779514508206e-21

* Branch 92
Rabr92 node_2 netRa92 319074756.9499282
Lbr92 netRa92 netL92 2.1786566800297914e-09
Rbbr92 netL92 0 -319115405.33306897
Cbr92 netL92 0 2.139691128491329e-26

* Branch 93
Rabr93 node_2 netRa93 -29416.29733412901
Lbr93 netRa93 netL93 -3.878229943785349e-11
Rbbr93 netL93 0 81287.83167631482
Cbr93 netL93 0 -1.624064374775514e-20

* Branch 94
Rabr94 node_2 netRa94 -48860.56899385352
Lbr94 netRa94 netL94 -2.8304846731745775e-11
Rbbr94 netL94 0 95390.00092669777
Cbr94 netL94 0 -6.077155442107245e-21

* Branch 95
Rabr95 node_2 netRa95 19716.38430100135
Lbr95 netRa95 netL95 -2.005535910616449e-11
Rbbr95 netL95 0 -83808.31207829215
Cbr95 netL95 0 -1.2117984041305945e-20

* Branch 96
Rabr96 node_2 netRa96 252070.6315270837
Lbr96 netRa96 netL96 1.0489128362495683e-10
Rbbr96 netL96 0 -407549.0243033612
Cbr96 netL96 0 1.021970182257888e-21

* Branch 97
Rabr97 node_2 netRa97 40003.868418291604
Lbr97 netRa97 netL97 3.503965345076338e-11
Rbbr97 netL97 0 -93199.0406174139
Cbr97 netL97 0 9.515931982677798e-21

* Branch 98
Rabr98 node_2 netRa98 -115521.52036047791
Lbr98 netRa98 netL98 3.899705358479186e-11
Rbbr98 netL98 0 133207.0511823642
Cbr98 netL98 0 2.493912306713945e-21

* Branch 99
Rabr99 node_2 netRa99 -59445.60805193387
Lbr99 netRa99 netL99 3.882227398017452e-11
Rbbr99 netL99 0 114931.9409793675
Cbr99 netL99 0 5.48462965582048e-21

.ends


.end
