* netlist generated with vector fitting poles and residues

.subckt total_network node_1 node_2 node_3 node_4 
X_11 node_1 0 yp11
X_12 node_1 node_2 yp12
X_13 node_1 node_3 yp13
X_14 node_1 node_4 yp14
X_22 node_2 0 yp22
X_23 node_2 node_3 yp23
X_24 node_2 node_4 yp24
X_33 node_3 0 yp33
X_34 node_3 node_4 yp34
X_44 node_4 0 yp44
.ends


* Y'11
.subckt yp11 node_1 0
* Branch 0
Rabr0 node_1 netRa0 1588.840361486932
Lbr0 netRa0 netL0 -9.817460440431366e-13
Rbbr0 netL0 0 -1982.7623076428276
Cbr0 netL0 0 -2.1614562516429894e-19

* Branch 1
Rabr1 node_1 netRa1 -1633200055925.8022
Lbr1 netRa1 netL1 0.0016921532282805148
Rbbr1 netL1 0 3918433649715.5425
Cbr1 netL1 0 2.642969830868501e-28

* Branch 2
Rabr2 node_1 netRa2 -361695825.900395
Lbr2 netRa2 netL2 -7.294402135094228e-07
Rbbr2 netL2 0 2400114052.5445685
Cbr2 netL2 0 -8.880196209578691e-25

* Branch 3
Rabr3 node_1 netRa3 49370367.98012091
Lbr3 netRa3 netL3 3.475009328287844e-08
Rbbr3 netL3 0 -82540065.65354721
Cbr3 netL3 0 8.81522444178443e-24

* Branch 4
Rabr4 node_1 netRa4 -58142268.58650153
Lbr4 netRa4 netL4 -4.1509660600371834e-09
Rbbr4 netL4 0 58533836.65686512
Cbr4 netL4 0 -1.2265893815421074e-24

* Branch 5
Rabr5 node_1 netRa5 2602616.279358712
Lbr5 netRa5 netL5 -5.15361650764126e-10
Rbbr5 netL5 0 -2734370.606270652
Cbr5 netL5 0 -7.108887986904487e-23

* Branch 6
Rabr6 node_1 netRa6 -983515499684.1316
Lbr6 netRa6 netL6 0.00029122303885330904
Rbbr6 netL6 0 1097004004204.2605
Cbr6 netL6 0 2.6940228191694637e-28

* Branch 7
Rabr7 node_1 netRa7 455.3923225649629
Lbr7 netRa7 netL7 1.627661400495288e-13
Rbbr7 netL7 0 -549.1187288079536
Cbr7 netL7 0 7.597769373193587e-19

* Branch 8
Rabr8 node_1 netRa8 3157.4081057929347
Lbr8 netRa8 netL8 -1.6182668752316053e-12
Rbbr8 netL8 0 -4245.061642168867
Cbr8 netL8 0 -1.1121985590224774e-19

* Branch 9
Rabr9 node_1 netRa9 -612.961246858263
Lbr9 netRa9 netL9 9.193837903837263e-13
Rbbr9 netL9 0 2455.5367072716695
Cbr9 netL9 0 5.396700876181662e-19

* Branch 10
Rabr10 node_1 netRa10 369905002211.9041
Lbr10 netRa10 netL10 0.00028024993001445097
Rbbr10 netL10 0 -693510131257.5963
Cbr10 netL10 0 1.0950107934495993e-27

* Branch 11
Rabr11 node_1 netRa11 21845.26361543776
Lbr11 netRa11 netL11 8.279999196310014e-12
Rbbr11 netL11 0 -26745.67841500572
Cbr11 netL11 0 1.448249067809507e-20

* Branch 12
Rabr12 node_1 netRa12 3880497.4349327423
Lbr12 netRa12 netL12 -3.4890896823746237e-10
Rbbr12 netL12 0 -3928286.877815363
Cbr12 netL12 0 -2.27885593076116e-23

* Branch 13
Rabr13 node_1 netRa13 -15928.707804035303
Lbr13 netRa13 netL13 -7.698507278705273e-12
Rbbr13 netL13 0 21776.967655182107
Cbr13 netL13 0 -2.2796682607212095e-20

* Branch 14
Rabr14 node_1 netRa14 39088.45401122913
Lbr14 netRa14 netL14 -4.8412862154671995e-12
Rbbr14 netL14 0 -39997.44215205381
Cbr14 netL14 0 -3.0559388255671234e-21

* Branch 15
Rabr15 node_1 netRa15 -31222083596856.41
Lbr15 netRa15 netL15 -0.007535405654486992
Rbbr15 netL15 0 34070614152673.43
Cbr15 netL15 0 -7.084495240842088e-30

* Branch 16
Rabr16 node_1 netRa16 -29.696703525330044
Lbr16 netRa16 netL16 6.259859954723005e-14
Rbbr16 netL16 0 156.3069045618295
Cbr16 netL16 0 8.066226109041928e-18

* Branch 17
Rabr17 node_1 netRa17 -203.16391756747498
Lbr17 netRa17 netL17 -2.9009615581749384e-13
Rbbr17 netL17 0 1181.164851236834
Cbr17 netL17 0 -1.7007568339566197e-18

* Branch 18
Rabr18 node_1 netRa18 5.501376061348831
Lbr18 netRa18 netL18 1.1433956320260308e-14
Rbbr18 netL18 0 40.20981032434526
Cbr18 netL18 0 5.1634495511472825e-17

* Branch 19
Rabr19 node_1 netRa19 1.8225791889849075
Lbr19 netRa19 netL19 2.6922249728504876e-12
Rbbr19 netL19 0 1014073.4889495556
Cbr19 netL19 0 2.163959372351222e-19

* Branch 20
Rabr20 node_1 netRa20 -73079343.88236074
Lbr20 netRa20 netL20 -2.1006264426027274e-07
Rbbr20 netL20 0 1183791865.909805
Cbr20 netL20 0 -2.532841684112728e-24

* Branch 21
Rabr21 node_1 netRa21 1181367.155508114
Lbr21 netRa21 netL21 2.9011443108519614e-09
Rbbr21 netL21 0 -14430850.84281968
Cbr21 netL21 0 1.7944823672951116e-22

* Branch 22
Rabr22 node_1 netRa22 -1109362.2958557042
Lbr22 netRa22 netL22 -2.7055387875690518e-09
Rbbr22 netL22 0 13394756.906048702
Cbr22 netL22 0 -1.9222009965815772e-22

* Branch 23
Rabr23 node_1 netRa23 3.2027794101539633
Lbr23 netRa23 netL23 1.1545404542090642e-13
Rbbr23 netL23 0 4714.1701826790795
Cbr23 netL23 0 4.9081794238671224e-18

* Branch 24
Rabr24 node_1 netRa24 -33657.485128589324
Lbr24 netRa24 netL24 -7.182513967734098e-12
Rbbr24 netL24 0 36530.193913261995
Cbr24 netL24 0 -6.068509489252549e-21

* Branch 25
Rd node_1 0 1838.4572499490437

.ends


* Y'12
.subckt yp12 node_1 node_2
* Branch 0
Rabr0 node_1 netRa0 -14068.43539754961
Lbr0 netRa0 netL0 -9.304314050411397e-12
Rbbr0 netL0 node_2 24997.74901951016
Cbr0 netL0 node_2 -5.018959733943971e-20

* Branch 1
Rabr1 node_1 netRa1 74161155274458.77
Lbr1 netRa1 netL1 -0.017549931689633525
Rbbr1 netL1 node_2 -79576372736030.73
Cbr1 netL1 node_2 -2.9735149208894263e-30

* Branch 2
Rabr2 node_1 netRa2 17.703186392976495
Lbr2 netRa2 netL2 8.585270876361667e-13
Rbbr2 netL2 node_2 186132.41080249316
Cbr2 netL2 node_2 8.884605551909033e-19

* Branch 3
Rabr3 node_1 netRa3 -28366765.82751658
Lbr3 netRa3 netL3 4.4973731865746195e-08
Rbbr3 netL3 node_2 115501569.98109034
Cbr3 netL3 node_2 1.2786671012982102e-23

* Branch 4
Rabr4 node_1 netRa4 174806.59996312266
Lbr4 netRa4 netL4 -1.1775336871760282e-09
Rbbr4 netL4 node_2 -6983910.341683773
Cbr4 netL4 node_2 -6.301820938527847e-22

* Branch 5
Rabr5 node_1 netRa5 50000.35223918096
Lbr5 netRa5 netL5 4.6249260076516934e-10
Rbbr5 netL5 node_2 -44402879.42801376
Cbr5 netL5 node_2 1.6421474614622508e-21

* Branch 6
Rabr6 node_1 netRa6 -131429183557.85854
Lbr6 netRa6 netL6 0.00027183557784627284
Rbbr6 netL6 node_2 862968952803.0259
Cbr6 netL6 node_2 2.3649382855061296e-27

* Branch 7
Rabr7 node_1 netRa7 -1017.6879622160087
Lbr7 netRa7 netL7 -1.521593365197246e-12
Rbbr7 netL7 node_2 8857.297206321968
Cbr7 netL7 node_2 -4.214529083312141e-19

* Branch 8
Rabr8 node_1 netRa8 221.32882769141412
Lbr8 netRa8 netL8 1.3181384201617715e-12
Rbbr8 netL8 node_2 -1920386.5168827167
Cbr8 netL8 node_2 5.328620881136727e-19

* Branch 9
Rabr9 node_1 netRa9 20923.011926781743
Lbr9 netRa9 netL9 5.971922281009161e-11
Rbbr9 netL9 node_2 -365051.2601712685
Cbr9 netL9 node_2 1.0437552233836552e-20

* Branch 10
Rabr10 node_1 netRa10 -1525512713452.752
Lbr10 netRa10 netL10 0.002363021712524802
Rbbr10 netL10 node_2 7064732249774.921
Cbr10 netL10 node_2 2.182159469670759e-28

* Branch 11
Rabr11 node_1 netRa11 234649.78249290877
Lbr11 netRa11 netL11 3.2086404175588697e-10
Rbbr11 netL11 node_2 -961313.2795924791
Cbr11 netL11 node_2 1.5418484232660048e-21

* Branch 12
Rabr12 node_1 netRa12 15234679.934157517
Lbr12 netRa12 netL12 6.504019796338935e-09
Rbbr12 netL12 node_2 -19573678.832981754
Cbr12 netL12 node_2 2.2275910200087237e-23

* Branch 13
Rabr13 node_1 netRa13 -194792.8770631409
Lbr13 netRa13 netL13 -3.4441954373918476e-10
Rbbr13 netL13 node_2 1226503.0007430615
Cbr13 netL13 node_2 -1.5960636706638729e-21

* Branch 14
Rabr14 node_1 netRa14 -8.491589289533332
Lbr14 netRa14 netL14 8.915870861173793e-13
Rbbr14 netL14 node_2 11728.435466181554
Cbr14 netL14 node_2 7.296273358350909e-19

* Branch 15
Rabr15 node_1 netRa15 -3893959015186.1577
Lbr15 netRa15 netL15 -0.009077301124596898
Rbbr15 netL15 node_2 37066123992272.36
Cbr15 netL15 node_2 -6.295272429730258e-29

* Branch 16
Rabr16 node_1 netRa16 -37.89989333047979
Lbr16 netRa16 netL16 2.9972213986139217e-13
Rbbr16 netL16 node_2 1117.9027300299117
Cbr16 netL16 node_2 2.0093080684865258e-18

* Branch 17
Rabr17 node_1 netRa17 101388.24601634826
Lbr17 netRa17 netL17 -1.0624802189010133e-11
Rbbr17 netL17 node_2 -103217.93473927146
Cbr17 netL17 node_2 -9.941608052009754e-22

* Branch 18
Rabr18 node_1 netRa18 77.93564789171523
Lbr18 netRa18 netL18 1.644920192451594e-13
Rbbr18 netL18 node_2 569.7964534187556
Cbr18 netL18 node_2 3.5890279936629765e-18

* Branch 19
Rabr19 node_1 netRa19 6011415308537.74
Lbr19 netRa19 netL19 -0.0043840182234510215
Rbbr19 netL19 node_2 -11478473831688.76
Cbr19 netL19 node_2 -6.329317680923964e-29

* Branch 20
Rabr20 node_1 netRa20 -6375052710.259946
Lbr20 netRa20 netL20 1.2039357704376986e-05
Rbbr20 netL20 node_2 45410380778.705765
Cbr20 netL20 node_2 4.0488336009144687e-26

* Branch 21
Rabr21 node_1 netRa21 31475353.8177509
Lbr21 netRa21 netL21 -1.7573063120273364e-07
Rbbr21 netL21 node_2 -1579844808.6277227
Cbr21 netL21 node_2 -3.162381127465992e-24

* Branch 22
Rabr22 node_1 netRa22 -25539712.71796491
Lbr22 netRa22 netL22 1.655655762062364e-07
Rbbr22 netL22 node_2 1685506302.50032
Cbr22 netL22 node_2 3.372851414868836e-24

* Branch 23
Rabr23 node_1 netRa23 -15999272.321992582
Lbr23 netRa23 netL23 -1.7164778940770292e-08
Rbbr23 netL23 node_2 51198262.12075853
Cbr23 netL23 node_2 -2.268148022261358e-23

* Branch 24
Rabr24 node_1 netRa24 934.5380909616373
Lbr24 netRa24 netL24 2.6477643253611056e-12
Rbbr24 netL24 node_2 -27794.372513480816
Cbr24 netL24 node_2 2.0229540613574216e-19

* Branch 25
Rd node_1 node_2 53018.326062394895

.ends


* Y'13
.subckt yp13 node_1 node_3
* Branch 0
Rabr0 node_1 netRa0 -6634.9007291937105
Lbr0 netRa0 netL0 -6.939710806081463e-12
Rbbr0 netL0 node_3 33584.34480914789
Cbr0 netL0 node_3 -1.2350303924859217e-19

* Branch 1
Rabr1 node_1 netRa1 -3262213362977.5947
Lbr1 netRa1 netL1 -0.002081228607439432
Rbbr1 netL1 node_3 4994157599702.44
Cbr1 netL1 node_3 -1.2778081833110277e-28

* Branch 2
Rabr2 node_1 netRa2 14.161990425516494
Lbr2 netRa2 netL2 6.868351767832106e-13
Rbbr2 netL2 node_3 148878.84458915738
Cbr2 netL2 node_3 1.110553869466212e-18

* Branch 3
Rabr3 node_1 netRa3 340427.25546139077
Lbr3 netRa3 netL3 5.710793712460595e-09
Rbbr3 netL3 node_3 -565792911.5994338
Cbr3 netL3 node_3 1.333996798842029e-22

* Branch 4
Rabr4 node_1 netRa4 -87601.00371205887
Lbr4 netRa4 netL4 -3.633250445795655e-10
Rbbr4 netL4 node_3 3027985.9651291533
Cbr4 netL4 node_3 -2.0342442780119218e-21

* Branch 5
Rabr5 node_1 netRa5 75882.00794839786
Lbr5 netRa5 netL5 1.8595487956714806e-10
Rbbr5 netL5 node_3 -855582.0232627867
Cbr5 netL5 node_3 3.726186368579456e-21

* Branch 6
Rabr6 node_1 netRa6 250514989228.00375
Lbr6 netRa6 netL6 7.104362295816299e-05
Rbbr6 netL6 node_3 -277130475298.8284
Cbr6 netL6 node_3 1.0251994241964171e-27

* Branch 7
Rabr7 node_1 netRa7 -536.1921800971659
Lbr7 netRa7 netL7 -1.2188419332413087e-12
Rbbr7 netL7 node_3 43698.986250922724
Cbr7 netL7 node_3 -5.871448597133283e-19

* Branch 8
Rabr8 node_1 netRa8 207.87538779425716
Lbr8 netRa8 netL8 1.0590993696238103e-12
Rbbr8 netL8 node_3 -51589.85142990035
Cbr8 netL8 node_3 6.605956550873131e-19

* Branch 9
Rabr9 node_1 netRa9 9792.18122127231
Lbr9 netRa9 netL9 3.678166734458526e-11
Rbbr9 netL9 node_3 -321744.5550493039
Cbr9 netL9 node_3 1.7429784347746746e-20

* Branch 10
Rabr10 node_1 netRa10 4062325426314.5337
Lbr10 netRa10 netL10 0.0015601336752910312
Rbbr10 netL10 node_3 -4974467019101.268
Cbr10 netL10 node_3 7.72956794198985e-29

* Branch 11
Rabr11 node_1 netRa11 202918.62213452876
Lbr11 netRa11 netL11 1.3557684805533073e-10
Rbbr11 netL11 node_3 -346767.6041611847
Cbr11 netL11 node_3 2.0025209571341002e-21

* Branch 12
Rabr12 node_1 netRa12 274169363.00934994
Lbr12 netRa12 netL12 1.2950610892887783e-08
Rbbr12 netL12 node_3 -275107497.976968
Cbr12 netL12 node_3 1.7209683086731272e-25

* Branch 13
Rabr13 node_1 netRa13 -191002.15152747594
Lbr13 netRa13 netL13 -1.386977394459019e-10
Rbbr13 netL13 node_3 351498.4091273382
Cbr13 netL13 node_3 -2.1513996121473328e-21

* Branch 14
Rabr14 node_1 netRa14 -3.307177371647908
Lbr14 netRa14 netL14 7.182399568205706e-13
Rbbr14 netL14 node_3 9859.530740419952
Cbr14 netL14 node_3 9.060750154985517e-19

* Branch 15
Rabr15 node_1 netRa15 -22797597061399.848
Lbr15 netRa15 netL15 -0.010018455611304954
Rbbr15 netL15 node_3 29693929567564.492
Cbr15 netL15 node_3 -1.4802135305835908e-29

* Branch 16
Rabr16 node_1 netRa16 -47.20022011388888
Lbr16 netRa16 netL16 2.4768475584281164e-13
Rbbr16 netL16 node_3 827.3406789626299
Cbr16 netL16 node_3 2.3731960580387126e-18

* Branch 17
Rabr17 node_1 netRa17 133597.37632095182
Lbr17 netRa17 netL17 -1.0722832031842813e-11
Rbbr17 netL17 node_3 -135018.59959327875
Cbr17 netL17 node_3 -5.849444870131297e-22

* Branch 18
Rabr18 node_1 netRa18 57.81829175276884
Lbr18 netRa18 netL18 1.3024429347160608e-13
Rbbr18 netL18 node_3 425.52522245164613
Cbr18 netL18 node_3 4.5291622833730164e-18

* Branch 19
Rabr19 node_1 netRa19 -63135383849663.29
Lbr19 netRa19 netL19 0.006050414479650887
Rbbr19 netL19 node_3 64130147656565.75
Cbr19 netL19 node_3 1.4935930350298112e-30

* Branch 20
Rabr20 node_1 netRa20 -5313743389.477623
Lbr20 netRa20 netL20 -5.444464667426045e-06
Rbbr20 netL20 node_3 15298197908.124935
Cbr20 netL20 node_3 -6.797660034248523e-26

* Branch 21
Rabr21 node_1 netRa21 107101797.61555876
Lbr21 netRa21 netL21 1.1593290482551484e-07
Rbbr21 netL21 node_3 -333578415.46699345
Cbr21 netL21 node_3 3.3206279746409434e-24

* Branch 22
Rabr22 node_1 netRa22 -103781130.25782944
Lbr22 netRa22 netL22 -1.1259846756193521e-07
Rbbr22 netL22 node_3 324413401.6239746
Cbr22 netL22 node_3 -3.424806644953065e-24

* Branch 23
Rabr23 node_1 netRa23 -32504070.180798635
Lbr23 netRa23 netL23 -2.8947048754232365e-08
Rbbr23 netL23 node_3 81098524.35416679
Cbr23 netL23 node_3 -1.1722064107649438e-23

* Branch 24
Rabr24 node_1 netRa24 784.4506910329702
Lbr24 netRa24 netL24 2.1214049127207605e-12
Rbbr24 netL24 node_3 -20444.793139430745
Cbr24 netL24 node_3 2.512486153314257e-19

* Branch 25
Rd node_1 node_3 28067.4605469162

.ends


* Y'14
.subckt yp14 node_1 node_4
* Branch 0
Rabr0 node_1 netRa0 -11945.683540315718
Lbr0 netRa0 netL0 -8.289766520709089e-12
Rbbr0 netL0 node_4 22635.75467532108
Cbr0 netL0 node_4 -6.084843390183328e-20

* Branch 1
Rabr1 node_1 netRa1 -14226093629938.975
Lbr1 netRa1 netL1 0.008667401924621506
Rbbr1 netL1 node_4 21110450743957.8
Cbr1 netL1 node_4 2.8852984219241703e-29

* Branch 2
Rabr2 node_1 netRa2 15.93278167740242
Lbr2 netRa2 netL2 7.726763712257281e-13
Rbbr2 netL2 node_4 167515.04241584582
Cbr2 netL2 node_4 9.871758510138295e-19

* Branch 3
Rabr3 node_1 netRa3 -7841908.497164179
Lbr3 netRa3 netL3 2.4902381902977332e-08
Rbbr3 netL3 node_4 98269034.20430844
Cbr3 netL3 node_4 2.8167856237455154e-23

* Branch 4
Rabr4 node_1 netRa4 56606.97806214401
Lbr4 netRa4 netL4 -9.1231910586263e-10
Rbbr4 netL4 node_4 -8569265.571590792
Cbr4 netL4 node_4 -8.287488662125749e-22

* Branch 5
Rabr5 node_1 netRa5 60351.40714177364
Lbr5 netRa5 netL5 3.796226122678576e-10
Rbbr5 netL5 node_4 -7791426.186977981
Cbr5 netL5 node_4 1.9873625423130285e-21

* Branch 6
Rabr6 node_1 netRa6 457431721537.8213
Lbr6 netRa6 netL6 0.0003067374107805956
Rbbr6 netL6 node_4 -729840362681.5519
Cbr6 netL6 node_4 9.22804266561051e-28

* Branch 7
Rabr7 node_1 netRa7 -888.3143361637354
Lbr7 netRa7 netL7 -1.3722551336706486e-12
Rbbr7 netL7 node_4 8575.183955867098
Cbr7 netL7 node_4 -4.732881900811365e-19

* Branch 8
Rabr8 node_1 netRa8 201.97316322820086
Lbr8 netRa8 netL8 1.186624615686574e-12
Rbbr8 netL8 node_4 -515962.92464868905
Cbr8 netL8 node_4 5.917557773660045e-19

* Branch 9
Rabr9 node_1 netRa9 18278.47188918518
Lbr9 netRa9 netL9 5.291343934562778e-11
Rbbr9 netL9 node_4 -329008.4306178066
Cbr9 netL9 node_4 1.1802022728442522e-20

* Branch 10
Rabr10 node_1 netRa10 19056273181368.465
Lbr10 netRa10 netL10 0.00627107665232574
Rbbr10 netL10 node_4 -22197403077018.254
Cbr10 netL10 node_4 1.4840309038992636e-29

* Branch 11
Rabr11 node_1 netRa11 228099.60724225687
Lbr11 netRa11 netL11 2.8385211656706613e-10
Rbbr11 netL11 node_4 -808736.2227183194
Cbr11 netL11 node_4 1.6553876660982102e-21

* Branch 12
Rabr12 node_1 netRa12 17502747.737685654
Lbr12 netRa12 netL12 6.3646139123011506e-09
Rbbr12 netL12 node_4 -21107928.259358514
Cbr12 netL12 node_4 1.75391916578654e-23

* Branch 13
Rabr13 node_1 netRa13 -194754.16337497853
Lbr13 netRa13 netL13 -3.0436956011417787e-10
Rbbr13 netL13 node_4 990732.9806639259
Cbr13 netL13 node_4 -1.7250138870018023e-21

* Branch 14
Rabr14 node_1 netRa14 -7.373391680797586
Lbr14 netRa14 netL14 8.026985706451477e-13
Rbbr14 netL14 node_4 10589.516170469285
Cbr14 netL14 node_4 8.10446640100217e-19

* Branch 15
Rabr15 node_1 netRa15 -1573813831988.714
Lbr15 netRa15 netL15 -0.012681468691937859
Rbbr15 netL15 node_4 162152012639350.03
Cbr15 netL15 node_4 -4.9861956342199145e-29

* Branch 16
Rabr16 node_1 netRa16 -35.59684197189401
Lbr16 netRa16 netL16 2.7082644276324354e-13
Rbbr16 netL16 node_4 1000.6662840794947
Cbr16 netL16 node_4 2.219845276422845e-18

* Branch 17
Rabr17 node_1 netRa17 96346.10347235911
Lbr17 netRa17 netL17 -9.817674834661025e-12
Rbbr17 netL17 node_4 -97991.06414970539
Cbr17 netL17 node_4 -1.018863130317038e-21

* Branch 18
Rabr18 node_1 netRa18 69.51040795339841
Lbr18 netRa18 netL18 1.479108687680583e-13
Rbbr18 netL18 node_4 508.38136323274904
Cbr18 netL18 node_4 3.9911936454212394e-18

* Branch 19
Rabr19 node_1 netRa19 2933883064611.9277
Lbr19 netRa19 netL19 -0.0027730224662853454
Rbbr19 netL19 node_4 -7410615452875.883
Cbr19 netL19 node_4 -1.269150538983755e-28

* Branch 20
Rabr20 node_1 netRa20 17476281792.07044
Lbr20 netRa20 netL20 9.954086917734008e-06
Rbbr20 netL20 node_4 -27557065453.338966
Cbr20 netL20 node_4 2.083965163078765e-26

* Branch 21
Rabr21 node_1 netRa21 -223776724.871803
Lbr21 netRa21 netL21 -1.701115830933298e-07
Rbbr21 netL21 node_4 455545915.86043507
Cbr21 netL21 node_4 -1.6958645891101486e-24

* Branch 22
Rabr22 node_1 netRa22 207918558.60056043
Lbr22 netRa22 netL22 1.6150305159195944e-07
Rbbr22 netL22 node_4 -432945173.185119
Cbr22 netL22 node_4 1.8248137292677318e-24

* Branch 23
Rabr23 node_1 netRa23 -17728404.456251938
Lbr23 netRa23 netL23 -1.65127008472062e-08
Rbbr23 netL23 node_4 46810697.66519667
Cbr23 netL23 node_4 -2.1305908135658613e-23

* Branch 24
Rabr24 node_1 netRa24 844.036932888092
Lbr24 netRa24 netL24 2.381463577963417e-12
Rbbr24 netL24 node_4 -24804.95056085302
Cbr24 netL24 node_4 2.248225936966883e-19

* Branch 25
Rd node_1 node_4 44392.92179200704

.ends


* Y'22
.subckt yp22 node_2 0
* Branch 0
Rabr0 node_2 netRa0 -58954.9558628037
Lbr0 netRa0 netL0 1.6865539133039877e-11
Rbbr0 netL0 0 62705.14503506671
Cbr0 netL0 0 3.7875280461454245e-21

* Branch 1
Rabr1 node_2 netRa1 483262683909.3987
Lbr1 netRa1 netL1 -0.0004079618013921675
Rbbr1 netL1 0 -932196764424.4861
Cbr1 netL1 0 -9.052515435278656e-28

* Branch 2
Rabr2 node_2 netRa2 -422286353.50089
Lbr2 netRa2 netL2 -2.788027494866112e-07
Rbbr2 netL2 0 667955541.3663424
Cbr2 netL2 0 -1.0061365597052839e-24

* Branch 3
Rabr3 node_2 netRa3 1.7267074159154696
Lbr3 netRa3 netL3 1.0874517039056703e-13
Rbbr3 netL3 0 4678.116691847138
Cbr3 netL3 0 7.012339555398884e-18

* Branch 4
Rabr4 node_2 netRa4 11902.52135724014
Lbr4 netRa4 netL4 1.0821476526610429e-10
Rbbr4 netL4 0 -4564987.969075276
Cbr4 netL4 0 7.015001129758108e-21

* Branch 5
Rabr5 node_2 netRa5 -2104.543255870554
Lbr5 netRa5 netL5 -4.037946058469483e-11
Rbbr5 netL5 0 -1254068.8083602197
Cbr5 netL5 0 -1.8861401368798793e-20

* Branch 6
Rabr6 node_2 netRa6 4776490279.797529
Lbr6 netRa6 netL6 4.658963281598257e-05
Rbbr6 netL6 0 -644557351224.8192
Cbr6 netL6 0 1.6157111771920026e-26

* Branch 7
Rabr7 node_2 netRa7 103.23561301683054
Lbr7 netRa7 netL7 9.159684806685169e-14
Rbbr7 netL7 0 -277.34306766184085
Cbr7 netL7 0 4.965625748861989e-18

* Branch 8
Rabr8 node_2 netRa8 33160.56808377571
Lbr8 netRa8 netL8 -7.187057007599652e-12
Rbbr8 netL8 0 -35300.59396079343
Cbr8 netL8 0 -5.925320137146321e-21

* Branch 9
Rabr9 node_2 netRa9 -221724.55017716013
Lbr9 netRa9 netL9 4.379346428836171e-11
Rbbr9 netL9 0 234582.8260692926
Cbr9 netL9 0 8.276058687485399e-22

* Branch 10
Rabr10 node_2 netRa10 -1850326089.0015397
Lbr10 netRa10 netL10 0.00019229051701497
Rbbr10 netL10 0 23012623500166.36
Cbr10 netL10 0 3.419861660273222e-27

* Branch 11
Rabr11 node_2 netRa11 -6801.998626431266
Lbr11 netRa11 netL11 2.5867579266606513e-12
Rbbr11 netL11 0 8273.384397789534
Cbr11 netL11 0 4.4996826816556e-20

* Branch 12
Rabr12 node_2 netRa12 -7340.094422244029
Lbr12 netRa12 netL12 -2.287365038154897e-11
Rbbr12 netL12 0 136000.28874291808
Cbr12 netL12 0 -2.7031436464345014e-20

* Branch 13
Rabr13 node_2 netRa13 14.173223964200242
Lbr13 netRa13 netL13 1.0697617798590694e-13
Rbbr13 netL13 0 -2119.4108128624152
Cbr13 netL13 0 6.068031337549072e-18

* Branch 14
Rabr14 node_2 netRa14 806517.9238289982
Lbr14 netRa14 netL14 5.7948028587109156e-11
Rbbr14 netL14 0 -812963.2679806205
Cbr14 netL14 0 8.906681846891534e-23

* Branch 15
Rabr15 node_2 netRa15 -621044528762.2833
Lbr15 netRa15 netL15 -0.000995216529676081
Rbbr15 netL15 0 3120416091539.3154
Cbr15 netL15 0 -5.138961500170224e-28

* Branch 16
Rabr16 node_2 netRa16 -1.149477422677617
Lbr16 netRa16 netL16 1.2392874065239952e-14
Rbbr16 netL16 0 49.4621125594789
Cbr16 netL16 0 4.9131554072253316e-17

* Branch 17
Rabr17 node_2 netRa17 -619266.7094114971
Lbr17 netRa17 netL17 -2.5983299441779366e-11
Rbbr17 netL17 0 621111.9880235317
Cbr17 netL17 0 -6.813232071937483e-23

* Branch 18
Rabr18 node_2 netRa18 170.82099815267557
Lbr18 netRa18 netL18 6.208214464596785e-13
Rbbr18 netL18 0 1567.627086680432
Cbr18 netL18 0 9.276801287634855e-19

* Branch 19
Rabr19 node_2 netRa19 -59660790715.48573
Lbr19 netRa19 netL19 -0.00024388825015724742
Rbbr19 netL19 0 1808404506561.0247
Cbr19 netL19 0 -2.3099329777989587e-27

* Branch 20
Rabr20 node_2 netRa20 0.7181994413781386
Lbr20 netRa20 netL20 1.116090377594092e-13
Rbbr20 netL20 0 24780.826338423536
Cbr20 netL20 0 5.080936639188462e-18

* Branch 21
Rabr21 node_2 netRa21 -922688.8810056222
Lbr21 netRa21 netL21 2.133379030578735e-09
Rbbr21 netL21 0 9218219.434929827
Cbr21 netL21 0 2.3918316799684167e-22

* Branch 22
Rabr22 node_2 netRa22 913802.5990853634
Lbr22 netRa22 netL22 -2.241355656779112e-09
Rbbr22 netL22 0 -10120522.725250933
Cbr22 netL22 0 -2.3013862260272925e-22

* Branch 23
Rabr23 node_2 netRa23 -9409187.625717673
Lbr23 netRa23 netL23 1.5714202414159383e-08
Rbbr23 netL23 0 50843332.83747555
Cbr23 netL23 0 2.936747839127317e-23

* Branch 24
Rabr24 node_2 netRa24 -6367937.805834998
Lbr24 netRa24 netL24 -3.438592972988886e-10
Rbbr24 netL24 0 6401757.505578161
Cbr24 netL24 0 -8.515470457986275e-24

* Branch 25
Rd node_2 0 10396.863933151462

.ends


* Y'23
.subckt yp23 node_2 node_3
* Branch 0
Rabr0 node_2 netRa0 -11154.341076757235
Lbr0 netRa0 netL0 -6.617139978262059e-12
Rbbr0 netL0 node_3 17536.735324056604
Cbr0 netL0 node_3 -5.874496448426861e-20

* Branch 1
Rabr1 node_2 netRa1 79697723411459.75
Lbr1 netRa1 netL1 -0.014271660291020626
Rbbr1 netL1 node_3 -83030110791538.27
Cbr1 netL1 node_3 -2.156548125114916e-30

* Branch 2
Rabr2 node_2 netRa2 12.392423847599932
Lbr2 netRa2 netL2 6.009649577955204e-13
Rbbr2 netL2 node_3 130301.71387584148
Cbr2 netL2 node_3 1.2692378135199123e-18

* Branch 3
Rabr3 node_2 netRa3 -45993498.450139515
Lbr3 netRa3 netL3 -3.7903643370825196e-08
Rbbr3 netL3 node_3 88599559.1208226
Cbr3 netL3 node_3 -9.671002805422863e-24

* Branch 4
Rabr4 node_2 netRa4 1850094.4456934296
Lbr4 netRa4 netL4 -1.886746239892106e-09
Rbbr4 netL4 node_3 -4190178.0077474327
Cbr4 netL4 node_3 -2.252856364088592e-22

* Branch 5
Rabr5 node_2 netRa5 -111126.84488573423
Lbr5 netRa5 netL5 4.998537741585192e-10
Rbbr5 netL5 node_3 2186844.154319466
Cbr5 netL5 node_3 1.4438220071725894e-21

* Branch 6
Rabr6 node_2 netRa6 -3688761229375.618
Lbr6 netRa6 netL6 -0.00041345750811004026
Rbbr6 netL6 node_3 3749913754175.932
Cbr6 netL6 node_3 -2.9912008064041656e-29

* Branch 7
Rabr7 node_2 netRa7 -793.7393415500842
Lbr7 netRa7 netL7 -1.0654077909841416e-12
Rbbr7 netL7 node_3 5067.602071370148
Cbr7 netL7 node_3 -5.735306846471599e-19

* Branch 8
Rabr8 node_2 netRa8 145.36807372036105
Lbr8 netRa8 netL8 9.212619614937578e-13
Rbbr8 netL8 node_3 143331.80791451872
Cbr8 netL8 node_3 7.632784462209701e-19

* Branch 9
Rabr9 node_2 netRa9 19306.09647562921
Lbr9 netRa9 netL9 4.733628519207893e-11
Rbbr9 netL9 node_3 -243061.677401842
Cbr9 netL9 node_3 1.2859069692358589e-20

* Branch 10
Rabr10 node_2 netRa10 -51887902701739.77
Lbr10 netRa10 netL10 -0.011886944319796679
Rbbr10 netL10 node_3 56031522965452.195
Cbr10 netL10 node_3 -4.09146291579318e-30

* Branch 11
Rabr11 node_2 netRa11 -80178.63093086208
Lbr11 netRa11 netL11 4.173890125321567e-10
Rbbr11 netL11 node_3 2644196.3165125283
Cbr11 netL11 node_3 1.5204797343933494e-21

* Branch 12
Rabr12 node_2 netRa12 -1885430.414451768
Lbr12 netRa12 netL12 4.7674948110123005e-09
Rbbr12 netL12 node_3 18300978.506165843
Cbr12 netL12 node_3 1.2296770817453022e-22

* Branch 13
Rabr13 node_2 netRa13 301852.2784551724
Lbr13 netRa13 netL13 -4.923449364588014e-10
Rbbr13 netL13 node_3 -1429980.6187008095
Cbr13 netL13 node_3 -1.0471473666068293e-21

* Branch 14
Rabr14 node_2 netRa14 -7.141535668153124
Lbr14 netRa14 netL14 6.224093370002863e-13
Rbbr14 netL14 node_3 8054.457146878078
Cbr14 netL14 node_3 1.0450042985348658e-18

* Branch 15
Rabr15 node_2 netRa15 -2032819019484.2263
Lbr15 netRa15 netL15 -0.004514869550489241
Rbbr15 netL15 node_3 17751758918142.7
Cbr15 netL15 node_3 -1.2523083747394896e-28

* Branch 16
Rabr16 node_2 netRa16 -21.74058086568606
Lbr16 netRa16 netL16 2.0776961362456142e-13
Rbbr16 netL16 node_3 808.9770151405053
Cbr16 netL16 node_3 2.9196543815097176e-18

* Branch 17
Rabr17 node_2 netRa17 61906.793677225774
Lbr17 netRa17 netL17 -6.994956391560974e-12
Rbbr17 netL17 node_3 -63203.522681786744
Cbr17 netL17 node_3 -1.7477462264867764e-21

* Branch 18
Rabr18 node_2 netRa18 55.75989154518441
Lbr18 netRa18 netL18 1.155473127650917e-13
Rbbr18 netL18 node_3 407.55425223965096
Cbr18 netL18 node_3 5.10947499561189e-18

* Branch 19
Rabr19 node_2 netRa19 2017845201603.1204
Lbr19 netRa19 netL19 -0.0015281242240272738
Rbbr19 netL19 node_3 -3996416827942.6226
Cbr19 netL19 node_3 -1.887478477418807e-28

* Branch 20
Rabr20 node_2 netRa20 -1778333041.939536
Lbr20 netRa20 netL20 3.6258368910910787e-06
Rbbr20 netL20 node_3 14443916314.373703
Cbr20 netL20 node_3 1.3713948813593349e-25

* Branch 21
Rabr21 node_2 netRa21 3760505.7713460266
Lbr21 netRa21 netL21 -6.26424251648998e-08
Rbbr21 netL21 node_3 -1366360410.3456209
Cbr21 netL21 node_3 -9.02684597130296e-24

* Branch 22
Rabr22 node_2 netRa22 -1897710.4945260019
Lbr22 netRa22 netL22 5.972404346907352e-08
Rbbr22 netL22 node_3 1973628587.0568275
Cbr22 netL22 node_3 9.484868094658577e-24

* Branch 23
Rabr23 node_2 netRa23 -10043619.058386989
Lbr23 netRa23 netL23 -1.0268720351674938e-08
Rbbr23 netL23 node_3 30033827.271218654
Cbr23 netL23 node_3 -3.670497566051581e-23

* Branch 24
Rabr24 node_2 netRa24 642.2425021041159
Lbr24 netRa24 netL24 1.8507392693785188e-12
Rbbr24 netL24 node_3 -20064.83715683441
Cbr24 netL24 node_3 2.8989802520605396e-19

* Branch 25
Rd node_2 node_3 42801.188061654844

.ends


* Y'24
.subckt yp24 node_2 node_4
* Branch 0
Rabr0 node_2 netRa0 -8468.317694429023
Lbr0 netRa0 netL0 -5.538901813270933e-12
Rbbr0 netL0 node_4 14839.917368792348
Cbr0 netL0 node_4 -8.279410566139621e-20

* Branch 1
Rabr1 node_2 netRa1 11735180362344.65
Lbr1 netRa1 netL1 -0.0035346970182367162
Rbbr1 netL1 node_4 -13123354523990.652
Cbr1 netL1 node_4 -2.2948837557394828e-29

* Branch 2
Rabr2 node_2 netRa2 10.621842153911274
Lbr2 netRa2 netL2 5.151150536837342e-13
Rbbr2 netL2 node_4 111677.57450584043
Cbr2 netL2 node_4 1.480771039815183e-18

* Branch 3
Rabr3 node_2 netRa3 -131860919.89031099
Lbr3 netRa3 netL3 7.786695370746728e-08
Rbbr3 netL3 node_4 190575696.42262512
Cbr3 netL3 node_4 3.016055701419818e-24

* Branch 4
Rabr4 node_2 netRa4 188167.2292018706
Lbr4 netRa4 netL4 -9.001560102940734e-10
Rbbr4 netL4 node_4 -4297555.981462035
Cbr4 netL4 node_4 -8.085111307198041e-22

* Branch 5
Rabr5 node_2 netRa5 27942.8994074866
Lbr5 netRa5 netL5 3.2353831953070323e-10
Rbbr5 netL5 node_4 52965794.5539746
Cbr5 netL5 node_4 2.351308385487309e-21

* Branch 6
Rabr6 node_2 netRa6 -1004328111032.8738
Lbr6 netRa6 netL6 0.00033603061748269943
Rbbr6 netL6 node_4 1152257788411.6882
Cbr6 netL6 node_4 2.897411281184429e-28

* Branch 7
Rabr7 node_2 netRa7 -625.201490250655
Lbr7 netRa7 netL7 -9.096141865252212e-13
Rbbr7 netL7 node_4 5009.074544553965
Cbr7 netL7 node_4 -6.9710422033352805e-19

* Branch 8
Rabr8 node_2 netRa8 129.957669591848
Lbr8 netRa8 netL8 7.910498854453346e-13
Rbbr8 netL8 node_4 425155.1374008171
Cbr8 netL8 node_4 8.882899659031001e-19

* Branch 9
Rabr9 node_2 netRa9 14504.08131296946
Lbr9 netRa9 netL9 3.77245202468831e-11
Rbbr9 netL9 node_4 -206881.23639391788
Cbr9 netL9 node_4 1.629877658776695e-20

* Branch 10
Rabr10 node_2 netRa10 638547866428.0476
Lbr10 netRa10 netL10 0.004860715884106654
Rbbr10 netL10 node_4 -58251807788402.734
Cbr10 netL10 node_4 1.3381787569714517e-28

* Branch 11
Rabr11 node_2 netRa11 131546.01161369568
Lbr11 netRa11 netL11 2.615045593590559e-10
Rbbr11 netL11 node_4 -1026618.9786384614
Cbr11 netL11 node_4 2.182047572917148e-21

* Branch 12
Rabr12 node_2 netRa12 5804222.036441839
Lbr12 netRa12 netL12 4.704570987271696e-09
Rbbr12 netL12 node_4 -11879325.558486745
Cbr12 netL12 node_4 7.104640438630606e-23

* Branch 13
Rabr13 node_2 netRa13 -77871.329752704
Lbr13 netRa13 netL13 -2.9062759024261624e-10
Rbbr13 netL13 node_4 2163718.0377902193
Cbr13 netL13 node_4 -2.1676731800442624e-21

* Branch 14
Rabr14 node_2 netRa14 -5.6227241995643995
Lbr14 netRa14 netL14 5.34382904824551e-13
Rbbr14 netL14 node_4 6970.63535467867
Cbr14 netL14 node_4 1.2172405285748423e-18

* Branch 15
Rabr15 node_2 netRa15 -344871036491.34973
Lbr15 netRa15 netL15 -0.003492488228084263
Rbbr15 netL15 node_4 55972903975318.92
Cbr15 netL15 node_4 -1.8170025720138552e-28

* Branch 16
Rabr16 node_2 netRa16 -21.4590163905655
Lbr16 netRa16 netL16 1.7926040334313073e-13
Rbbr16 netL16 node_4 677.3281031369869
Cbr16 netL16 node_4 3.3672717773784944e-18

* Branch 17
Rabr17 node_2 netRa17 58092.429072905536
Lbr17 netRa17 netL17 -6.245770686524613e-12
Rbbr17 netL17 node_4 -59195.34225735302
Cbr17 netL17 node_4 -1.7775556309382856e-21

* Branch 18
Rabr18 node_2 netRa18 46.962681022593635
Lbr18 netRa18 netL18 9.8770620988249e-14
Rbbr18 netL18 node_4 343.3113623786424
Cbr18 netL18 node_4 5.9772263829630625e-18

* Branch 19
Rabr19 node_2 netRa19 485648650896.8197
Lbr19 netRa19 netL19 -0.0009417065773017672
Rbbr19 netL19 node_4 -3588520714567.5713
Cbr19 netL19 node_4 -5.349244867843851e-28

* Branch 20
Rabr20 node_2 netRa20 286216451.48023885
Lbr20 netRa20 netL20 4.003436093301739e-06
Rbbr20 netL20 node_4 -123894619046.47798
Cbr20 netL20 node_4 1.413166083220085e-25

* Branch 21
Rabr21 node_2 netRa21 -18336605.72526114
Lbr21 netRa21 netL21 -7.188955140101395e-08
Rbbr21 netL21 node_4 560100981.7818589
Cbr21 netL21 node_4 -7.629214887721211e-24

* Branch 22
Rabr22 node_2 netRa22 18456758.726673834
Lbr22 netRa22 netL22 6.856436065728759e-08
Rbbr22 netL22 node_4 -506938747.7677256
Cbr22 netL22 node_4 7.968799963390935e-24

* Branch 23
Rabr23 node_2 netRa23 -9755791.240585454
Lbr23 netRa23 netL23 -9.761016338104757e-09
Rbbr23 netL23 node_4 28319987.912952866
Cbr23 netL23 node_4 -3.8029681290187584e-23

* Branch 24
Rabr24 node_2 netRa24 557.0257125294409
Lbr24 netRa24 netL24 1.5873518811746534e-12
Rbbr24 netL24 node_4 -16846.382978754013
Cbr24 netL24 node_4 3.376314996466647e-19

* Branch 25
Rd node_2 node_4 32154.700991568145

.ends


* Y'33
.subckt yp33 node_3 0
* Branch 0
Rabr0 node_3 netRa0 -869.0439590030843
Lbr0 netRa0 netL0 -2.201184519943969e-12
Rbbr0 netL0 0 -5567.62079883981
Cbr0 netL0 0 -5.609716050955061e-19

* Branch 1
Rabr1 node_3 netRa1 -7732611212317012.0
Lbr1 netRa1 netL1 -0.08586607568945336
Rbbr1 netL1 0 7733854596566434.0
Cbr1 netL1 0 -1.435825077268484e-33

* Branch 2
Rabr2 node_3 netRa2 284600040.6260958
Lbr2 netRa2 netL2 4.541046616365462e-07
Rbbr2 netL2 0 -1276824924.7672884
Cbr2 netL2 0 1.305189742227765e-24

* Branch 3
Rabr3 node_3 netRa3 -10169646.055456707
Lbr3 netRa3 netL3 -1.4724738458886085e-08
Rbbr3 netL3 0 40151238.132258266
Cbr3 netL3 0 -3.865634647084155e-23

* Branch 4
Rabr4 node_3 netRa4 81613.60912161233
Lbr4 netRa4 netL4 1.1166512872792313e-10
Rbbr4 netL4 0 -306594.120314986
Cbr4 netL4 0 5.001630560318261e-21

* Branch 5
Rabr5 node_3 netRa5 4.924828640199055
Lbr5 netRa5 netL5 1.225413332314085e-13
Rbbr5 netL5 0 2968.2491779127863
Cbr5 netL5 0 6.215035733076237e-18

* Branch 6
Rabr6 node_3 netRa6 196304155201.06473
Lbr6 netRa6 netL6 -0.00010985794458169535
Rbbr6 netL6 0 -277078463737.8788
Cbr6 netL6 0 -2.0124372509579626e-27

* Branch 7
Rabr7 node_3 netRa7 625.6734779086544
Lbr7 netRa7 netL7 -5.114040221374794e-13
Rbbr7 netL7 0 -1060.203819476362
Cbr7 netL7 0 -5.806588710983281e-19

* Branch 8
Rabr8 node_3 netRa8 14240.673859258924
Lbr8 netRa8 netL8 9.157122374549406e-12
Rbbr8 netL8 0 -23630.911722735727
Cbr8 netL8 0 3.04833712241556e-20

* Branch 9
Rabr9 node_3 netRa9 -6042.710421662218
Lbr9 netRa9 netL9 -2.444994659148616e-11
Rbbr9 netL9 0 238251.45177771765
Cbr9 netL9 0 -2.6357937950120823e-20

* Branch 10
Rabr10 node_3 netRa10 715694960258.1718
Lbr10 netRa10 netL10 -0.0005560654453030678
Rbbr10 netL10 0 -1371059848216.4502
Cbr10 netL10 0 -5.653301857844264e-28

* Branch 11
Rabr11 node_3 netRa11 -616.0243659165337
Lbr11 netRa11 netL11 -2.4279718037857347e-12
Rbbr11 netL11 0 19439.145602498786
Cbr11 netL11 0 -2.6101481346581924e-19

* Branch 12
Rabr12 node_3 netRa12 2354065.024710437
Lbr12 netRa12 netL12 2.8732992883401885e-10
Rbbr12 netL12 0 -2408046.1650481075
Cbr12 netL12 0 5.0991361951483356e-23

* Branch 13
Rabr13 node_3 netRa13 2.8389946662685475
Lbr13 netRa13 netL13 1.1173666347256627e-13
Rbbr13 netL13 0 5827.687240432968
Cbr13 netL13 0 5.851466746682312e-18

* Branch 14
Rabr14 node_3 netRa14 654.1995523587844
Lbr14 netRa14 netL14 9.951760328013371e-12
Rbbr14 netL14 0 366847.6153737407
Cbr14 netL14 0 6.553198095344975e-20

* Branch 15
Rabr15 node_3 netRa15 -2531587757522.2363
Lbr15 netRa15 netL15 -0.0017661328400582464
Rbbr15 netL15 0 4461807095713.475
Cbr15 netL15 0 -1.5640374069978698e-28

* Branch 16
Rabr16 node_3 netRa16 0.4657054908605407
Lbr16 netRa16 netL16 1.640564097093815e-14
Rbbr16 netL16 0 90.17352453125459
Cbr16 netL16 0 3.8193409824396444e-17

* Branch 17
Rabr17 node_3 netRa17 -3127.9782661413687
Lbr17 netRa17 netL17 -1.824518657385588e-12
Rbbr17 netL17 0 5153.225742345985
Cbr17 netL17 0 -1.2835301281834039e-19

* Branch 18
Rabr18 node_3 netRa18 151.6201275555534
Lbr18 netRa18 netL18 1.57968865312354e-13
Rbbr18 netL18 0 101934.92555001147
Cbr18 netL18 0 3.2924561409865182e-18

* Branch 19
Rabr19 node_3 netRa19 201585313288.51376
Lbr19 netRa19 netL19 0.00024209027183394916
Rbbr19 netL19 0 -703782841680.1993
Cbr19 netL19 0 1.7171895189162406e-27

* Branch 20
Rabr20 node_3 netRa20 111210650.47466025
Lbr20 netRa20 netL20 -2.3103762865969346e-07
Rbbr20 netL20 0 -933087689.6767405
Cbr20 netL20 0 -2.1618831970335846e-24

* Branch 21
Rabr21 node_3 netRa21 2.23480417879234
Lbr21 netRa21 netL21 1.240349442489519e-13
Rbbr21 netL21 0 72230.61459852
Cbr21 netL21 0 4.571628081072184e-18

* Branch 22
Rabr22 node_3 netRa22 -102928.51183111989
Lbr22 netRa22 netL22 2.0755935638779173e-10
Rbbr22 netL22 0 810216.6540095113
Cbr22 netL22 0 2.384795722509077e-21

* Branch 23
Rabr23 node_3 netRa23 -246815.32532878552
Lbr23 netRa23 netL23 -1.8362430942783444e-09
Rbbr23 netL23 0 51349043.36872266
Cbr23 netL23 0 -3.069106305262124e-22

* Branch 24
Rabr24 node_3 netRa24 -87416.62078751018
Lbr24 netRa24 netL24 -2.6555285480682243e-11
Rbbr24 netL24 0 102788.51086873871
Cbr24 netL24 0 -3.1214085173285328e-21

* Branch 25
Rd node_3 0 3864.9781911711675

.ends


* Y'34
.subckt yp34 node_3 node_4
* Branch 0
Rabr0 node_3 netRa0 -14012.715082792969
Lbr0 netRa0 netL0 -9.986306295089626e-12
Rbbr0 netL0 node_4 27598.301836989725
Cbr0 netL0 node_4 -5.264986291820307e-20

* Branch 1
Rabr1 node_3 netRa1 -160712030353736.9
Lbr1 netRa1 netL1 0.03423950226023431
Rbbr1 netL1 node_4 170223606307008.9
Cbr1 netL1 node_4 1.2514659581092235e-30

* Branch 2
Rabr2 node_3 netRa2 19.473181704808955
Lbr2 netRa2 netL2 9.443820693986516e-13
Rbbr2 netL2 node_4 204732.87186965923
Cbr2 netL2 node_4 8.076894733262426e-19

* Branch 3
Rabr3 node_3 netRa3 -7449729.683137421
Lbr3 netRa3 netL3 3.196801340699465e-08
Rbbr3 netL3 node_4 157548826.37846723
Cbr3 netL3 node_4 2.2717466872135907e-23

* Branch 4
Rabr4 node_3 netRa4 482.3325376057071
Lbr4 netRa4 netL4 -1.1619499584222743e-09
Rbbr4 netL4 node_4 -19281776.8315135
Cbr4 netL4 node_4 -6.550128421368503e-22

* Branch 5
Rabr5 node_3 netRa5 100101.10996047758
Lbr5 netRa5 netL5 4.813173755683874e-10
Rbbr5 netL5 node_4 -5673690.037796682
Cbr5 netL5 node_4 1.5518296619373088e-21

* Branch 6
Rabr6 node_3 netRa6 566278100516.8757
Lbr6 netRa6 netL6 0.00027671423928491123
Rbbr6 netL6 node_4 -745145616610.9216
Cbr6 netL6 node_4 6.578731415177318e-28

* Branch 7
Rabr7 node_3 netRa7 -1073.062811301462
Lbr7 netRa7 netL7 -1.6692082552395433e-12
Rbbr7 netL7 node_4 10596.578972288846
Cbr7 netL7 node_4 -3.900996695700992e-19

* Branch 8
Rabr8 node_3 netRa8 246.0671264768681
Lbr8 netRa8 netL8 1.451714137213641e-12
Rbbr8 netL8 node_4 -804943.8340194474
Cbr8 netL8 node_4 4.837400100971458e-19

* Branch 9
Rabr9 node_3 netRa9 24926.10172739368
Lbr9 netRa9 netL9 6.592786017269303e-11
Rbbr9 netL9 node_4 -368532.89047854074
Cbr9 netL9 node_4 9.351102975956043e-21

* Branch 10
Rabr10 node_3 netRa10 12606389007851.027
Lbr10 netRa10 netL10 -0.004510006627595497
Rbbr10 netL10 node_4 -15057051138487.969
Cbr10 netL10 node_4 -2.3733820891713466e-29

* Branch 11
Rabr11 node_3 netRa11 415897.61087126733
Lbr11 netRa11 netL11 4.6146297665875696e-10
Rbbr11 netL11 node_4 -1250689.231291274
Cbr11 netL11 node_4 9.466427981923747e-22

* Branch 12
Rabr12 node_3 netRa12 51482576.693421505
Lbr12 netRa12 netL12 1.4745064167023348e-08
Rbbr12 netL12 node_4 -58035818.70878522
Cbr12 netL12 node_4 5.0051103370650564e-24

* Branch 13
Rabr13 node_3 netRa13 -351554.53617792914
Lbr13 netRa13 netL13 -5.079468221256191e-10
Rbbr13 netL13 node_4 1571031.6169845855
Cbr13 netL13 node_4 -9.986639940125342e-22

* Branch 14
Rabr14 node_3 netRa14 -9.744209099982914
Lbr14 netRa14 netL14 9.807976935146224e-13
Rbbr14 netL14 node_4 12857.19492901435
Cbr14 netL14 node_4 6.632400036354326e-19

* Branch 15
Rabr15 node_3 netRa15 -5804185548500.216
Lbr15 netRa15 netL15 -0.009276351166785548
Rbbr15 netL15 node_4 29038544590887.71
Cbr15 netL15 node_4 -5.507484693620786e-29

* Branch 16
Rabr16 node_3 netRa16 -43.30168292098268
Lbr16 netRa16 netL16 3.308215981253953e-13
Rbbr16 netL16 node_4 1223.592106986643
Cbr16 netL16 node_4 1.817618920366317e-18

* Branch 17
Rabr17 node_3 netRa17 116375.50770935169
Lbr17 netRa17 netL17 -1.1938299722754127e-11
Rbbr17 netL17 node_4 -118388.93888993878
Cbr17 netL17 node_4 -8.488650010076987e-22

* Branch 18
Rabr18 node_3 netRa18 84.73694244518354
Lbr18 netRa18 netL18 1.8072659639279625e-13
Rbbr18 netL18 node_4 619.8230941496237
Cbr18 netL18 node_4 3.2664362069325563e-18

* Branch 19
Rabr19 node_3 netRa19 5763590513537.1875
Lbr19 netRa19 netL19 -0.003834807931416363
Rbbr19 netL19 node_4 -10127991698054.389
Cbr19 netL19 node_4 -6.546623754249597e-29

* Branch 20
Rabr20 node_3 netRa20 2546253165.322754
Lbr20 netRa20 netL20 7.000489487532445e-06
Rbbr20 netL20 node_4 -37884073223.60219
Cbr20 netL20 node_4 7.555883206692294e-26

* Branch 21
Rabr21 node_3 netRa21 -81842136.78945255
Lbr21 netRa21 netL21 -1.3776927936177074e-07
Rbbr21 netL21 node_4 505867187.95343107
Cbr21 netL21 node_4 -3.449881108685571e-24

* Branch 22
Rabr22 node_3 netRa22 80452076.43347113
Lbr22 netRa22 netL22 1.322812925610312e-07
Rbbr22 netL22 node_4 -478192263.505021
Cbr22 netL22 node_4 3.565305805740242e-24

* Branch 23
Rabr23 node_3 netRa23 -21555948.577822816
Lbr23 netRa23 netL23 -1.959754490337117e-08
Rbbr23 netL23 node_4 55188804.218639426
Cbr23 netL23 node_4 -1.760944705517195e-23

* Branch 24
Rabr24 node_3 netRa24 1029.2510267127957
Lbr24 netRa24 netL24 2.9089789697509435e-12
Rbbr24 netL24 node_4 -30396.10752240365
Cbr24 netL24 node_4 1.840847436553574e-19

* Branch 25
Rd node_3 node_4 52605.313194775365

.ends


* Y'44
.subckt yp44 node_4 0
* Branch 0
Rabr0 node_4 netRa0 13137.987775185315
Lbr0 netRa0 netL0 -5.10699795382105e-12
Rbbr0 netL0 0 -14592.407869250419
Cbr0 netL0 0 -2.0845067672488893e-20

* Branch 1
Rabr1 node_4 netRa1 8092354615908.762
Lbr1 netRa1 netL1 0.004884418508311415
Rbbr1 netL1 0 -11937838783997.01
Cbr1 netL1 0 5.057387607380292e-29

* Branch 2
Rabr2 node_4 netRa2 -232938517.86843824
Lbr2 netRa2 netL2 2.625861460692296e-07
Rbbr2 netL2 0 609718900.9257227
Cbr2 netL2 0 1.794889287249321e-24

* Branch 3
Rabr3 node_4 netRa3 4775796.392075933
Lbr3 netRa3 netL3 -6.131728234491008e-09
Rbbr3 netL3 0 -14523360.874326104
Cbr3 netL3 0 -8.343701059819436e-23

* Branch 4
Rabr4 node_4 netRa4 4.071173924510055
Lbr4 netRa4 netL4 1.1989134154531737e-13
Rbbr4 netL4 0 3511.6056453241417
Cbr4 netL4 0 6.355701478947164e-18

* Branch 5
Rabr5 node_4 netRa5 -5318.258325157871
Lbr5 netRa5 netL5 1.9221999335385255e-11
Rbbr5 netL5 0 73447.62260109285
Cbr5 netL5 0 3.669140107069949e-20

* Branch 6
Rabr6 node_4 netRa6 1340802220145.1084
Lbr6 netRa6 netL6 0.00028998211948928033
Rbbr6 netL6 0 -1423616515309.8708
Cbr6 netL6 0 1.5213334399840861e-28

* Branch 7
Rabr7 node_4 netRa7 3318.872029927979
Lbr7 netRa7 netL7 -1.0397911877175245e-12
Rbbr7 netL7 0 -3718.317581920918
Cbr7 netL7 0 -7.485476291764152e-20

* Branch 8
Rabr8 node_4 netRa8 3762.399662474082
Lbr8 netRa8 netL8 3.783354034750926e-12
Rbbr8 netL8 0 -10270.708067733192
Cbr8 netL8 0 1.1765669734659758e-19

* Branch 9
Rabr9 node_4 netRa9 -85006.63527717932
Lbr9 netRa9 netL9 -2.9123349855592425e-11
Rbbr9 netL9 0 100565.0009827536
Cbr9 netL9 0 -3.51254683156314e-21

* Branch 10
Rabr10 node_4 netRa10 171309482280.0506
Lbr10 netRa10 netL10 -0.0001887791446721607
Rbbr10 netL10 0 -486557153830.4719
Cbr10 netL10 0 -2.2571755507055383e-27

* Branch 11
Rabr11 node_4 netRa11 -8348.731020976238
Lbr11 netRa11 netL11 5.620208861522673e-12
Rbbr11 netL11 0 13917.264096492872
Cbr11 netL11 0 4.6593872564903307e-20

* Branch 12
Rabr12 node_4 netRa12 1.6629156401676823
Lbr12 netRa12 netL12 1.1234744482413235e-13
Rbbr12 netL12 0 5041.910219536679
Cbr12 netL12 0 5.819427290804645e-18

* Branch 13
Rabr13 node_4 netRa13 3817.8331032207916
Lbr13 netRa13 netL13 -3.704726876254078e-12
Rbbr13 netL13 0 -9041.460467705272
Cbr13 netL13 0 -1.0191223522576653e-19

* Branch 14
Rabr14 node_4 netRa14 9628.050568420886
Lbr14 netRa14 netL14 8.265739923339178e-12
Rbbr14 netL14 0 -21634.928542353755
Cbr14 netL14 0 4.3709145089404277e-20

* Branch 15
Rabr15 node_4 netRa15 -171580609934.50748
Lbr15 netRa15 netL15 -0.0013120801948070158
Rbbr15 netL15 0 15936002419454.156
Cbr15 netL15 0 -4.814075632118243e-28

* Branch 16
Rabr16 node_4 netRa16 0.4248607324322415
Lbr16 netRa16 netL16 1.559031337783043e-14
Rbbr16 netL16 0 85.37429642367056
Cbr16 netL16 0 4.018329191145346e-17

* Branch 17
Rabr17 node_4 netRa17 -7046.367318568103
Lbr17 netRa17 netL17 -2.5674553089808842e-12
Rbbr17 netL17 0 8741.407335549495
Cbr17 netL17 0 -4.5004003398148336e-20

* Branch 18
Rabr18 node_4 netRa18 122.24709570466999
Lbr18 netRa18 netL18 1.8302213561399853e-13
Rbbr18 netL18 0 1072.9818118539142
Cbr18 netL18 0 3.1608297750262943e-18

* Branch 19
Rabr19 node_4 netRa19 9947779945909.676
Lbr19 netRa19 netL19 0.0015780480119030689
Rbbr19 netL19 0 -10377826352645.463
Cbr19 netL19 0 1.529848348087236e-29

* Branch 20
Rabr20 node_4 netRa20 266011741.1986874
Lbr20 netRa20 netL20 -2.3566483831020986e-07
Rbbr20 netL20 0 -629559560.768326
Cbr20 netL20 0 -1.3895061947121537e-24

* Branch 21
Rabr21 node_4 netRa21 -116217.14175956002
Lbr21 netRa21 netL21 2.6827038030943724e-10
Rbbr21 netL21 0 1157746.7002141248
Cbr21 netL21 0 1.9014584226786004e-21

* Branch 22
Rabr22 node_4 netRa22 2.196000523503705
Lbr22 netRa22 netL22 1.2057046366536008e-13
Rbbr22 netL22 0 61958.10427957007
Cbr22 netL22 0 4.702975861278944e-18

* Branch 23
Rabr23 node_4 netRa23 -1364074.5506347024
Lbr23 netRa23 netL23 -2.647041941598082e-09
Rbbr23 netL23 0 11883465.629899496
Cbr23 netL23 0 -1.8937440988076625e-22

* Branch 24
Rabr24 node_4 netRa24 -329895.2444511353
Lbr24 netRa24 netL24 -5.3551918503371256e-11
Rbbr24 netL24 0 346038.03128666244
Cbr24 netL24 0 -4.828347678171704e-22

* Branch 25
Rd node_4 0 2904.2777211518032

.ends


.end
