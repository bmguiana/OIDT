* netlist generated with vector fitting poles and residues

.subckt total_network node_1 node_2 node_3 node_4 
X_11 node_1 0 yp11
X_12 node_1 node_2 yp12
X_13 node_1 node_3 yp13
X_14 node_1 node_4 yp14
X_22 node_2 0 yp22
X_23 node_2 node_3 yp23
X_24 node_2 node_4 yp24
X_33 node_3 0 yp33
X_34 node_3 node_4 yp34
X_44 node_4 0 yp44
.ends


* Y'11
.subckt yp11 node_1 0
* Branch 0
Rabr0 node_1 netRa0 9682.55713555277
Lbr0 netRa0 netL0 -1.3057374482872816e-11
Rbbr0 netL0 0 -65093.07268096887
Cbr0 netL0 0 -2.0005385540770708e-20

* Branch 1
Rabr1 node_1 netRa1 -114.34416309868016
Lbr1 netRa1 netL1 -2.8677797070629378e-11
Rbbr1 netL1 0 -4207687.046794687
Cbr1 netL1 0 -1.3041157784312053e-20

* Branch 2
Rabr2 node_1 netRa2 10450.205590163956
Lbr2 netRa2 netL2 -1.43591505855453e-11
Rbbr2 netL2 0 -73197.99111794688
Cbr2 netL2 0 -1.823535239063292e-20

* Branch 3
Rabr3 node_1 netRa3 14830.563171383776
Lbr3 netRa3 netL3 -2.21778197117018e-11
Rbbr3 netL3 0 -106086.9536937453
Cbr3 netL3 0 -1.3672189493273814e-20

* Branch 4
Rabr4 node_1 netRa4 45685.540439772056
Lbr4 netRa4 netL4 -5.944952230663264e-11
Rbbr4 netL4 0 -168767.93110950515
Cbr4 netL4 0 -7.521869188143886e-21

* Branch 5
Rabr5 node_1 netRa5 -46444.88689428135
Lbr5 netRa5 netL5 -4.555961872515317e-11
Rbbr5 netL5 0 162958.53448667488
Cbr5 netL5 0 -6.1341594638928334e-21

* Branch 6
Rabr6 node_1 netRa6 756458.5129565139
Lbr6 netRa6 netL6 2.2158946513337628e-10
Rbbr6 netL6 0 -866715.7803845919
Cbr6 netL6 0 3.3986499359415727e-22

* Branch 7
Rabr7 node_1 netRa7 992315.8271891995
Lbr7 netRa7 netL7 1.8409278134796681e-10
Rbbr7 netL7 0 -1077372.5147544127
Cbr7 netL7 0 1.7279675873309792e-22

* Branch 8
Rabr8 node_1 netRa8 -18832.469095122036
Lbr8 netRa8 netL8 -1.0223041711423415e-10
Rbbr8 netL8 0 920743.9500050528
Cbr8 netL8 0 -6.557244623371741e-21

* Branch 9
Rabr9 node_1 netRa9 51555.394195445566
Lbr9 netRa9 netL9 -4.8367070734926385e-11
Rbbr9 netL9 0 -156629.85828399024
Cbr9 netL9 0 -5.896467785420137e-21

* Branch 10
Rabr10 node_1 netRa10 11324.87518919889
Lbr10 netRa10 netL10 -9.71637947391237e-11
Rbbr10 netL10 0 -671272.4850327042
Cbr10 netL10 0 -1.1178575530008759e-20

* Branch 11
Rabr11 node_1 netRa11 41469.10900646528
Lbr11 netRa11 netL11 -6.480869518416271e-11
Rbbr11 netL11 0 -179418.17680649023
Cbr11 netL11 0 -8.499628905015623e-21

* Branch 12
Rabr12 node_1 netRa12 57134.12619653855
Lbr12 netRa12 netL12 -2.2280861615706043e-11
Rbbr12 netL12 0 -82588.70685229654
Cbr12 netL12 0 -4.693200724672375e-21

* Branch 13
Rabr13 node_1 netRa13 21259.937631155386
Lbr13 netRa13 netL13 -7.147655923838164e-11
Rbbr13 netL13 0 -304275.9791640061
Cbr13 netL13 0 -1.0496649020162748e-20

* Branch 14
Rabr14 node_1 netRa14 -22379.599743931645
Lbr14 netRa14 netL14 -2.2399993926125166e-11
Rbbr14 netL14 0 92040.82727598262
Cbr14 netL14 0 -1.1039095644377212e-20

* Branch 15
Rabr15 node_1 netRa15 3051.3690189883255
Lbr15 netRa15 netL15 -1.2214986870949049e-11
Rbbr15 netL15 0 -151373.20765029188
Cbr15 netL15 0 -2.5007529426912268e-20

* Branch 16
Rabr16 node_1 netRa16 56053.82667127487
Lbr16 netRa16 netL16 -4.272171391083969e-11
Rbbr16 netL16 0 -161807.68478213297
Cbr16 netL16 0 -4.6599189176663524e-21

* Branch 17
Rabr17 node_1 netRa17 16705.887340598456
Lbr17 netRa17 netL17 -7.765142569707275e-11
Rbbr17 netL17 0 -406829.4161683298
Cbr17 netL17 0 -1.0752226292840858e-20

* Branch 18
Rabr18 node_1 netRa18 -12621.372756057304
Lbr18 netRa18 netL18 -1.3177319270599409e-10
Rbbr18 netL18 0 2824601.6757770134
Cbr18 netL18 0 -4.285754795544353e-21

* Branch 19
Rabr19 node_1 netRa19 11435.619093261614
Lbr19 netRa19 netL19 -8.410376146685486e-11
Rbbr19 netL19 0 -600545.6984765135
Cbr19 netL19 0 -1.1187206478676762e-20

* Branch 20
Rabr20 node_1 netRa20 22870.25711686823
Lbr20 netRa20 netL20 -6.780817119144698e-11
Rbbr20 netL20 0 -279417.95244734123
Cbr20 netL20 0 -1.0232627403648788e-20

* Branch 21
Rabr21 node_1 netRa21 3665.4652504473356
Lbr21 netRa21 netL21 -1.0206972447223453e-10
Rbbr21 netL21 0 -1597373.5097560373
Cbr21 netL21 0 -1.2955689191095389e-20

* Branch 22
Rabr22 node_1 netRa22 11037704.4933524
Lbr22 netRa22 netL22 7.116321640066881e-10
Rbbr22 netL22 0 -11149588.967409648
Cbr22 netL22 0 5.78697233842848e-24

* Branch 23
Rabr23 node_1 netRa23 18715.46971047185
Lbr23 netRa23 netL23 -4.5030529344377164e-11
Rbbr23 netL23 0 -178918.0632834639
Cbr23 netL23 0 -1.3087705704887156e-20

* Branch 24
Rabr24 node_1 netRa24 7122.9953706235265
Lbr24 netRa24 netL24 -8.758918681358107e-11
Rbbr24 netL24 0 -948104.112885361
Cbr24 netL24 0 -1.138993802952057e-20

* Branch 25
Rabr25 node_1 netRa25 26246.24464171199
Lbr25 netRa25 netL25 -4.7403613239620146e-11
Rbbr25 netL25 0 -214955.11012955688
Cbr25 netL25 0 -8.235447948274391e-21

* Branch 26
Rabr26 node_1 netRa26 9131.850507255338
Lbr26 netRa26 netL26 -6.168011436586669e-11
Rbbr26 netL26 0 -776375.9563538962
Cbr26 netL26 0 -8.150117383381276e-21

* Branch 27
Rabr27 node_1 netRa27 1907.922450095985
Lbr27 netRa27 netL27 -8.56764015091066e-11
Rbbr27 netL27 0 -1645838.3127996193
Cbr27 netL27 0 -1.907436904283744e-20

* Branch 28
Rabr28 node_1 netRa28 25044555.436964214
Lbr28 netRa28 netL28 -1.4302322633121214e-09
Rbbr28 netL28 0 -25088582.543713357
Cbr28 netL28 0 -2.275014491614527e-24

* Branch 29
Rabr29 node_1 netRa29 11936.41441889433
Lbr29 netRa29 netL29 -8.996425243799957e-11
Rbbr29 netL29 0 -417093.8244735396
Cbr29 netL29 0 -1.6932037987337186e-20

* Branch 30
Rabr30 node_1 netRa30 -2039.812479780282
Lbr30 netRa30 netL30 -8.11547536647565e-11
Rbbr30 netL30 0 9038849.467473593
Cbr30 netL30 0 -6.704438981515437e-21

* Branch 31
Rabr31 node_1 netRa31 169169784.70056576
Lbr31 netRa31 netL31 -2.9161342194399864e-09
Rbbr31 netL31 0 -169249481.0021429
Cbr31 netL31 0 -1.0183544104148048e-25

* Branch 32
Rabr32 node_1 netRa32 17857.268611137908
Lbr32 netRa32 netL32 -7.88403086596318e-11
Rbbr32 netL32 0 -384571.915619451
Cbr32 netL32 0 -1.1099632005335666e-20

* Branch 33
Rabr33 node_1 netRa33 -2808.7776832747395
Lbr33 netRa33 netL33 -8.52374144298187e-11
Rbbr33 netL33 0 2309554.5937944558
Cbr33 netL33 0 -1.7097393641934817e-20

* Branch 34
Rabr34 node_1 netRa34 14984.735604828786
Lbr34 netRa34 netL34 -8.962831364910095e-11
Rbbr34 netL34 0 -264698.3010156331
Cbr34 netL34 0 -2.1611026381641544e-20

* Branch 35
Rabr35 node_1 netRa35 -65944.29758979697
Lbr35 netRa35 netL35 -1.970941125207198e-10
Rbbr35 netL35 0 401155.6924110156
Cbr35 netL35 0 -7.608958998679423e-21

* Branch 36
Rabr36 node_1 netRa36 233753.18454862852
Lbr36 netRa36 netL36 -1.6289096019701788e-10
Rbbr36 netL36 0 -328883.141154217
Cbr36 netL36 0 -2.1090352341135614e-21

* Branch 37
Rabr37 node_1 netRa37 248521.28326171817
Lbr37 netRa37 netL37 -2.0185016442036176e-10
Rbbr37 netL37 0 -354917.8402061073
Cbr37 netL37 0 -2.276671842672379e-21

* Branch 38
Rabr38 node_1 netRa38 163289.15597340005
Lbr38 netRa38 netL38 -1.2596535819630183e-10
Rbbr38 netL38 0 -312180.940634655
Cbr38 netL38 0 -2.459024596174798e-21

* Branch 39
Rabr39 node_1 netRa39 3921.8718088871656
Lbr39 netRa39 netL39 -6.8948072256909e-11
Rbbr39 netL39 0 -898096.0764479276
Cbr39 netL39 0 -1.7618068585068034e-20

* Branch 40
Rabr40 node_1 netRa40 26112.461428301165
Lbr40 netRa40 netL40 -3.6809835260050025e-11
Rbbr40 netL40 0 -180962.21770745743
Cbr40 netL40 0 -7.729413568700118e-21

* Branch 41
Rabr41 node_1 netRa41 23407.136065766197
Lbr41 netRa41 netL41 -4.6016342413184756e-11
Rbbr41 netL41 0 -224556.78643393956
Cbr41 netL41 0 -8.66288095453309e-21

* Branch 42
Rabr42 node_1 netRa42 -111817.41997280526
Lbr42 netRa42 netL42 -2.549220928717159e-10
Rbbr42 netL42 0 462439.507942023
Cbr42 netL42 0 -4.98680040192516e-21

* Branch 43
Rabr43 node_1 netRa43 115834.98793769428
Lbr43 netRa43 netL43 -1.7466881228158853e-10
Rbbr43 netL43 0 -450398.34694360686
Cbr43 netL43 0 -3.327747783277522e-21

* Branch 44
Rabr44 node_1 netRa44 4770113.481247232
Lbr44 netRa44 netL44 4.120651190001868e-10
Rbbr44 netL44 0 -4873610.1495759655
Cbr44 netL44 0 1.773112085312013e-23

* Branch 45
Rabr45 node_1 netRa45 -69585.12138403358
Lbr45 netRa45 netL45 -8.423099949188626e-11
Rbbr45 netL45 0 419518.74372744234
Cbr45 netL45 0 -2.8974229142809013e-21

* Branch 46
Rabr46 node_1 netRa46 -10079.371338638643
Lbr46 netRa46 netL46 -1.7121637089127173e-11
Rbbr46 netL46 0 112852.17369184022
Cbr46 netL46 0 -1.5136107145254464e-20

* Branch 47
Rabr47 node_1 netRa47 14565.286634803382
Lbr47 netRa47 netL47 -5.4140078834884714e-11
Rbbr47 netL47 0 -428102.0631348831
Cbr47 netL47 0 -8.582773221954248e-21

* Branch 48
Rabr48 node_1 netRa48 97229.26005092342
Lbr48 netRa48 netL48 -1.7846704880354776e-10
Rbbr48 netL48 0 -240906.12999013995
Cbr48 netL48 0 -7.577769813541472e-21

* Branch 49
Rabr49 node_1 netRa49 338767.1130435258
Lbr49 netRa49 netL49 -2.5347077327062853e-10
Rbbr49 netL49 0 -523208.1258627136
Cbr49 netL49 0 -1.4273545883037223e-21

* Branch 50
Rabr50 node_1 netRa50 46215.700704076706
Lbr50 netRa50 netL50 -1.0358516441408545e-10
Rbbr50 netL50 0 -390624.9462871416
Cbr50 netL50 0 -5.7065660438796865e-21

* Branch 51
Rabr51 node_1 netRa51 -204652.0137794727
Lbr51 netRa51 netL51 -4.096591572887711e-10
Rbbr51 netL51 0 672465.8948864035
Cbr51 netL51 0 -2.988719583426691e-21

* Branch 52
Rabr52 node_1 netRa52 46573.32753899094
Lbr52 netRa52 netL52 1.4512539540052528e-10
Rbbr52 netL52 0 -372108.89665791334
Cbr52 netL52 0 8.424927182135198e-21

* Branch 53
Rabr53 node_1 netRa53 1726536.3592950145
Lbr53 netRa53 netL53 -4.235817804260487e-10
Rbbr53 netL53 0 -2010074.856853814
Cbr53 netL53 0 -1.2200702036542217e-22

* Branch 54
Rabr54 node_1 netRa54 19238.253698783617
Lbr54 netRa54 netL54 -1.7825870372506728e-10
Rbbr54 netL54 0 -700173.7350087942
Cbr54 netL54 0 -1.3048272039136972e-20

* Branch 55
Rabr55 node_1 netRa55 -35161.98219027599
Lbr55 netRa55 netL55 -2.147567241326797e-10
Rbbr55 netL55 0 1101071.3639419975
Cbr55 netL55 0 -5.595027481463152e-21

* Branch 56
Rabr56 node_1 netRa56 -131737485.51209903
Lbr56 netRa56 netL56 1.0901180536805525e-09
Rbbr56 netL56 0 131765610.3056443
Cbr56 netL56 0 6.279963310308649e-26

* Branch 57
Rabr57 node_1 netRa57 77167849.80705222
Lbr57 netRa57 netL57 4.472308716672802e-09
Rbbr57 netL57 0 -77393865.78123914
Cbr57 netL57 0 7.488962250241873e-25

* Branch 58
Rabr58 node_1 netRa58 106519.9164418697
Lbr58 netRa58 netL58 -1.999366344823068e-10
Rbbr58 netL58 0 -1084093.1503970383
Cbr58 netL58 0 -1.727365077600453e-21

* Branch 59
Rabr59 node_1 netRa59 84783.97306374945
Lbr59 netRa59 netL59 -2.3945322339132947e-10
Rbbr59 netL59 0 -975618.450176162
Cbr59 netL59 0 -2.8859798055025494e-21

* Branch 60
Rabr60 node_1 netRa60 -274032.96352520015
Lbr60 netRa60 netL60 -2.638192846848659e-10
Rbbr60 netL60 0 540378.953311806
Cbr60 netL60 0 -1.7834301546492213e-21

* Branch 61
Rabr61 node_1 netRa61 154298.29042904548
Lbr61 netRa61 netL61 -3.428231761719265e-10
Rbbr61 netL61 0 -507961.6170379043
Cbr61 netL61 0 -4.3655152379207156e-21

* Branch 62
Rabr62 node_1 netRa62 86442.23437768547
Lbr62 netRa62 netL62 -1.8423978126581513e-10
Rbbr62 netL62 0 -1132671.0804320984
Cbr62 netL62 0 -1.8783032101037832e-21

* Branch 63
Rabr63 node_1 netRa63 94201.65807350216
Lbr63 netRa63 netL63 -1.9176923733257716e-10
Rbbr63 netL63 0 -1001998.1040704352
Cbr63 netL63 0 -2.0281888208235348e-21

* Branch 64
Rabr64 node_1 netRa64 114302.1183012913
Lbr64 netRa64 netL64 1.7280268638337392e-10
Rbbr64 netL64 0 -695094.0015162415
Cbr64 netL64 0 2.177372535309686e-21

* Branch 65
Rabr65 node_1 netRa65 354842.00570296723
Lbr65 netRa65 netL65 2.3341389959530434e-10
Rbbr65 netL65 0 -618691.9900351671
Cbr65 netL65 0 1.0637062146869933e-21

* Branch 66
Rabr66 node_1 netRa66 447302.1304621728
Lbr66 netRa66 netL66 -4.271915734254416e-10
Rbbr66 netL66 0 -920322.0276496577
Cbr66 netL66 0 -1.0370230968358913e-21

* Branch 67
Rabr67 node_1 netRa67 376558.38534929074
Lbr67 netRa67 netL67 -3.059346425704384e-10
Rbbr67 netL67 0 -655377.9794246895
Cbr67 netL67 0 -1.2389802211811195e-21

* Branch 68
Rabr68 node_1 netRa68 1085154.3630374959
Lbr68 netRa68 netL68 -3.901748552694756e-10
Rbbr68 netL68 0 -1374587.3995451198
Cbr68 netL68 0 -2.6151173737517833e-22

* Branch 69
Rabr69 node_1 netRa69 34548.60363424101
Lbr69 netRa69 netL69 -1.973003403894922e-10
Rbbr69 netL69 0 -1859974.5220063783
Cbr69 netL69 0 -3.0591283886078028e-21

* Branch 70
Rabr70 node_1 netRa70 -46610.82992682521
Lbr70 netRa70 netL70 -3.365338474005415e-10
Rbbr70 netL70 0 1934911.549437783
Cbr70 netL70 0 -3.747085174210252e-21

* Branch 71
Rabr71 node_1 netRa71 -66375.79126875788
Lbr71 netRa71 netL71 -1.7597250571783944e-10
Rbbr71 netL71 0 722504.0753517589
Cbr71 netL71 0 -3.674984968442499e-21

* Branch 72
Rabr72 node_1 netRa72 172197.43254405973
Lbr72 netRa72 netL72 -4.1564491171888284e-10
Rbbr72 netL72 0 -662888.5019494534
Cbr72 netL72 0 -3.636276997932023e-21

* Branch 73
Rabr73 node_1 netRa73 29347.96717728647
Lbr73 netRa73 netL73 -6.257884433755777e-10
Rbbr73 netL73 0 -9839112.626600254
Cbr73 netL73 0 -2.1450596104908287e-21

* Branch 74
Rabr74 node_1 netRa74 -11224.021294439988
Lbr74 netRa74 netL74 -2.9989431436463247e-10
Rbbr74 netL74 0 18457099.917889107
Cbr74 netL74 0 -1.4652635162234554e-21

* Branch 75
Rabr75 node_1 netRa75 -156486.37523366843
Lbr75 netRa75 netL75 2.47247881849154e-10
Rbbr75 netL75 0 982508.3701259521
Cbr75 netL75 0 1.6070777240820507e-21

* Branch 76
Rabr76 node_1 netRa76 -24084.209798688382
Lbr76 netRa76 netL76 -2.719888493101353e-10
Rbbr76 netL76 0 1242262.16152548
Cbr76 netL76 0 -9.129012673132862e-21

* Branch 77
Rabr77 node_1 netRa77 7937.0248223572125
Lbr77 netRa77 netL77 -2.6165644724500296e-10
Rbbr77 netL77 0 -11617045.454573656
Cbr77 netL77 0 -2.8048063029532962e-21

* Branch 78
Rabr78 node_1 netRa78 1121699.3974779765
Lbr78 netRa78 netL78 -8.828689188553905e-10
Rbbr78 netL78 0 -1595217.1237832112
Cbr78 netL78 0 -4.932679776459767e-22

* Branch 79
Rabr79 node_1 netRa79 -126839.59069689907
Lbr79 netRa79 netL79 -5.586772753253861e-10
Rbbr79 netL79 0 2617870.4561887933
Cbr79 netL79 0 -1.685044677051499e-21

* Branch 80
Rabr80 node_1 netRa80 1714023.837914427
Lbr80 netRa80 netL80 -5.896895323295918e-10
Rbbr80 netL80 0 -2101821.61759149
Cbr80 netL80 0 -1.6366881272818276e-22

* Branch 81
Rabr81 node_1 netRa81 14714808.150913727
Lbr81 netRa81 netL81 2.267725577194213e-09
Rbbr81 netL81 0 -15348371.668686816
Cbr81 netL81 0 1.0041269173146611e-23

* Branch 82
Rabr82 node_1 netRa82 2568512.6257469854
Lbr82 netRa82 netL82 -1.7322120941551782e-09
Rbbr82 netL82 0 -3625937.012569474
Cbr82 netL82 0 -1.8596791343269728e-22

* Branch 83
Rabr83 node_1 netRa83 382935.1538786665
Lbr83 netRa83 netL83 -1.0219753144397296e-09
Rbbr83 netL83 0 -2944651.663113624
Cbr83 netL83 0 -9.058961007313597e-22

* Branch 84
Rabr84 node_1 netRa84 12823012.574129483
Lbr84 netRa84 netL84 -2.6964125115956525e-09
Rbbr84 netL84 0 -13878403.10997521
Cbr84 netL84 0 -1.5151398752781792e-23

* Branch 85
Rabr85 node_1 netRa85 6234846.680932968
Lbr85 netRa85 netL85 -1.5556690571699668e-09
Rbbr85 netL85 0 -6995887.115323972
Cbr85 netL85 0 -3.566521953051848e-23

* Branch 86
Rabr86 node_1 netRa86 2470211.5844459627
Lbr86 netRa86 netL86 -9.048513350972868e-10
Rbbr86 netL86 0 -3188406.6928252876
Cbr86 netL86 0 -1.1488427410817078e-22

* Branch 87
Rabr87 node_1 netRa87 11534331.586890833
Lbr87 netRa87 netL87 -2.155225476930708e-09
Rbbr87 netL87 0 -12344267.435059767
Cbr87 netL87 0 -1.513666535250697e-23

* Branch 88
Rabr88 node_1 netRa88 1064670.4459916332
Lbr88 netRa88 netL88 -5.654332369364657e-10
Rbbr88 netL88 0 -1594733.7372524485
Cbr88 netL88 0 -3.3299769378386537e-22

* Branch 89
Rabr89 node_1 netRa89 7460827.359669573
Lbr89 netRa89 netL89 1.7198370574088764e-09
Rbbr89 netL89 0 -7936214.396692571
Cbr89 netL89 0 2.904738064759144e-23

* Branch 90
Rabr90 node_1 netRa90 294823.15503231314
Lbr90 netRa90 netL90 -3.94285706210743e-10
Rbbr90 netL90 0 -566359.0378465967
Cbr90 netL90 0 -2.360615299949183e-21

* Branch 91
Rabr91 node_1 netRa91 977994.6978583133
Lbr91 netRa91 netL91 6.495665551504662e-10
Rbbr91 netL91 0 -1512539.3067362758
Cbr91 netL91 0 4.391992619172064e-22

* Branch 92
Rabr92 node_1 netRa92 -384261.5760588635
Lbr92 netRa92 netL92 1.8247440383364183e-10
Rbbr92 netL92 0 605557.9405767513
Cbr92 netL92 0 7.840352380927874e-22

* Branch 93
Rabr93 node_1 netRa93 -762463.9093596427
Lbr93 netRa93 netL93 3.004728875957946e-10
Rbbr93 netL93 0 1044709.8522855884
Cbr93 netL93 0 3.771503517754213e-22

* Branch 94
Rabr94 node_1 netRa94 -179076.6149656584
Lbr94 netRa94 netL94 1.7834617836727172e-10
Rbbr94 netL94 0 674063.7839210406
Cbr94 netL94 0 1.4767312622198368e-21

* Branch 95
Rabr95 node_1 netRa95 -92652.8971422058
Lbr95 netRa95 netL95 1.232067406742945e-10
Rbbr95 netL95 0 558840.2636198879
Cbr95 netL95 0 2.3770251979808217e-21

* Branch 96
Rabr96 node_1 netRa96 -115088.91782996857
Lbr96 netRa96 netL96 3.9934131097917535e-11
Rbbr96 netL96 0 158936.1408476183
Cbr96 netL96 0 2.1823813989942028e-21

* Branch 97
Rabr97 node_1 netRa97 -209399.30955134015
Lbr97 netRa97 netL97 4.859909689596806e-11
Rbbr97 netL97 0 245797.732884778
Cbr97 netL97 0 9.439862907825367e-22

* Branch 98
Rabr98 node_1 netRa98 28404.64963254128
Lbr98 netRa98 netL98 4.0284223826521204e-11
Rbbr98 netL98 0 -228612.88879784456
Cbr98 netL98 0 6.227738761727498e-21

* Branch 99
Rabr99 node_1 netRa99 -5825.083924182491
Lbr99 netRa99 netL99 8.331465805279803e-12
Rbbr99 netL99 0 44561.489849757156
Cbr99 netL99 0 3.171759814695979e-20

.ends


* Y'12
.subckt yp12 node_1 node_2
* Branch 0
Rabr0 node_1 netRa0 -62.58069107566079
Lbr0 netRa0 netL0 -1.8539132900532938e-13
Rbbr0 netL0 node_2 990.6010491386801
Cbr0 netL0 node_2 -5.495423195913943e-18

* Branch 1
Rabr1 node_1 netRa1 -62.21373002579572
Lbr1 netRa1 netL1 -1.8924516320552873e-13
Rbbr1 netL1 node_2 857.942184449639
Cbr1 netL1 node_2 -5.5622872860030776e-18

* Branch 2
Rabr2 node_1 netRa2 -1432.6654811164756
Lbr2 netRa2 netL2 7.148274216489782e-13
Rbbr2 netL2 node_2 2408.335293632243
Cbr2 netL2 node_2 2.0051075476174338e-19

* Branch 3
Rabr3 node_1 netRa3 -514.3957072856632
Lbr3 netRa3 netL3 -6.452093867445039e-13
Rbbr3 netL3 node_2 2935.6654974148
Cbr3 netL3 node_2 -4.624696622565695e-19

* Branch 4
Rabr4 node_1 netRa4 -109375.48678455772
Lbr4 netRa4 netL4 1.52049275074209e-11
Rbbr4 netL4 node_2 115097.35253143254
Cbr4 netL4 node_2 1.1992185237017718e-21

* Branch 5
Rabr5 node_1 netRa5 -57.49044210952698
Lbr5 netRa5 netL5 -2.0871222846654754e-13
Rbbr5 netL5 node_2 692.2843452108765
Cbr5 netL5 node_2 -6.33620217535906e-18

* Branch 6
Rabr6 node_1 netRa6 1.4619523144589839
Lbr6 netRa6 netL6 -2.0616635294962343e-13
Rbbr6 netL6 node_2 -12045.115363304882
Cbr6 netL6 node_2 -1.7503027104604437e-18

* Branch 7
Rabr7 node_1 netRa7 -99.79776433344638
Lbr7 netRa7 netL7 7.152775890350326e-14
Rbbr7 netL7 node_2 245.91659604609933
Cbr7 netL7 node_2 2.8378420804851562e-18

* Branch 8
Rabr8 node_1 netRa8 -684.7549483044369
Lbr8 netRa8 netL8 -2.7355302919124925e-13
Rbbr8 netL8 node_2 990.0073740525363
Cbr8 netL8 node_2 -4.0955296706741242e-19

* Branch 9
Rabr9 node_1 netRa9 -954.8366093872069
Lbr9 netRa9 netL9 2.0273664994784765e-13
Rbbr9 netL9 node_2 1100.6273552537402
Cbr9 netL9 node_2 1.9144695584438997e-19

* Branch 10
Rabr10 node_1 netRa10 7610.802261489743
Lbr10 netRa10 netL10 -7.642501421187337e-13
Rbbr10 netL10 node_2 -7876.154083022356
Cbr10 netL10 node_2 -1.2705918402286374e-20

* Branch 11
Rabr11 node_1 netRa11 -152.18028438492564
Lbr11 netRa11 netL11 1.1750007471395472e-13
Rbbr11 netL11 node_2 453.47468860087724
Cbr11 netL11 node_2 1.661612761726029e-18

* Branch 12
Rabr12 node_1 netRa12 -57.286108972104316
Lbr12 netRa12 netL12 -2.0955380041693255e-13
Rbbr12 netL12 node_2 658.3783854983067
Cbr12 netL12 node_2 -6.227126331363145e-18

* Branch 13
Rabr13 node_1 netRa13 154.53183509261112
Lbr13 netRa13 netL13 1.1686054595652173e-13
Rbbr13 netL13 node_2 -460.3911337576766
Cbr13 netL13 node_2 1.6785384146039946e-18

* Branch 14
Rabr14 node_1 netRa14 -25.53013086880497
Lbr14 netRa14 netL14 -1.109845957339489e-13
Rbbr14 netL14 node_2 1125.0274337292553
Cbr14 netL14 node_2 -4.321343405461276e-18

* Branch 15
Rabr15 node_1 netRa15 -62.35345959017306
Lbr15 netRa15 netL15 -1.9213229913253063e-13
Rbbr15 netL15 node_2 627.2812527064984
Cbr15 netL15 node_2 -5.30861209800123e-18

* Branch 16
Rabr16 node_1 netRa16 -501.5870672620703
Lbr16 netRa16 netL16 3.6702819477697156e-13
Rbbr16 netL16 node_2 1375.1020217498913
Cbr16 netL16 node_2 5.233544991225334e-19

* Branch 17
Rabr17 node_1 netRa17 9.34321398793786
Lbr17 netRa17 netL17 -9.730555393331334e-14
Rbbr17 netL17 node_2 -1875.6076978748401
Cbr17 netL17 node_2 -4.524883459033538e-18

* Branch 18
Rabr18 node_1 netRa18 -9.804416504426209
Lbr18 netRa18 netL18 -1.0184274620869301e-13
Rbbr18 netL18 node_2 2971.560790255816
Cbr18 netL18 node_2 -4.47566264430685e-18

* Branch 19
Rabr19 node_1 netRa19 89289.96312225914
Lbr19 netRa19 netL19 -2.51290689451615e-12
Rbbr19 netL19 node_2 -89477.49603721466
Cbr19 netL19 node_2 -3.1435328920988226e-22

* Branch 20
Rabr20 node_1 netRa20 -59.42806265159106
Lbr20 netRa20 netL20 -2.0856819478048247e-13
Rbbr20 netL20 node_2 621.5809437400084
Cbr20 netL20 node_2 -6.016926082794956e-18

* Branch 21
Rabr21 node_1 netRa21 -48.21768523094178
Lbr21 netRa21 netL21 -1.2076476233302352e-13
Rbbr21 netL21 node_2 638.7414594894476
Cbr21 netL21 node_2 -4.093712896238499e-18

* Branch 22
Rabr22 node_1 netRa22 -53.92523418992264
Lbr22 netRa22 netL22 -2.1451257388759233e-13
Rbbr22 netL22 node_2 629.1301927330903
Cbr22 netL22 node_2 -6.772100285146472e-18

* Branch 23
Rabr23 node_1 netRa23 -30.19488435504372
Lbr23 netRa23 netL23 -1.4023659204673002e-13
Rbbr23 netL23 node_2 1192.8715796883303
Cbr23 netL23 node_2 -4.215927016099918e-18

* Branch 24
Rabr24 node_1 netRa24 -517.6498899928202
Lbr24 netRa24 netL24 -2.48640014706122e-13
Rbbr24 netL24 node_2 838.8826959954695
Cbr24 netL24 node_2 -5.771266452232396e-19

* Branch 25
Rabr25 node_1 netRa25 16.95649902719069
Lbr25 netRa25 netL25 4.403887672240018e-13
Rbbr25 netL25 node_2 -51482.65908422327
Cbr25 netL25 node_2 8.763388245216724e-19

* Branch 26
Rabr26 node_1 netRa26 -156.3234116283897
Lbr26 netRa26 netL26 8.989252726740378e-13
Rbbr26 netL26 node_2 15379.851953589005
Cbr26 netL26 node_2 3.4275898605164103e-19

* Branch 27
Rabr27 node_1 netRa27 -862.4588893182901
Lbr27 netRa27 netL27 -4.573656722669933e-13
Rbbr27 netL27 node_2 1552.5328060510942
Cbr27 netL27 node_2 -3.4394153981497186e-19

* Branch 28
Rabr28 node_1 netRa28 8.859689523074115
Lbr28 netRa28 netL28 -1.2537136254106608e-13
Rbbr28 netL28 node_2 -5115.743347749456
Cbr28 netL28 node_2 -2.3414118531002054e-18

* Branch 29
Rabr29 node_1 netRa29 -59.12158137443745
Lbr29 netRa29 netL29 -1.5785245957477006e-13
Rbbr29 netL29 node_2 630.5720562851552
Cbr29 netL29 node_2 -4.373046988161978e-18

* Branch 30
Rabr30 node_1 netRa30 -60.65600982191219
Lbr30 netRa30 netL30 -1.6026286647968268e-13
Rbbr30 netL30 node_2 587.9658450755225
Cbr30 netL30 node_2 -4.632348856590795e-18

* Branch 31
Rabr31 node_1 netRa31 -491.82534957397354
Lbr31 netRa31 netL31 -3.7678936214277116e-13
Rbbr31 netL31 node_2 1331.7974888781744
Cbr31 netL31 node_2 -5.802272309208809e-19

* Branch 32
Rabr32 node_1 netRa32 -23.45235047222287
Lbr32 netRa32 netL32 -1.3472022712012963e-13
Rbbr32 netL32 node_2 1273.1180144435411
Cbr32 netL32 node_2 -4.792808596512668e-18

* Branch 33
Rabr33 node_1 netRa33 100.02014718170315
Lbr33 netRa33 netL33 -1.475150144933886e-13
Rbbr33 netL33 node_2 -619.3657081296749
Cbr33 netL33 node_2 -2.34723131588011e-18

* Branch 34
Rabr34 node_1 netRa34 -64.85600243436076
Lbr34 netRa34 netL34 -1.7648170651437114e-13
Rbbr34 netL34 node_2 587.6853205718126
Cbr34 netL34 node_2 -4.756384406866584e-18

* Branch 35
Rabr35 node_1 netRa35 -55.032020035601924
Lbr35 netRa35 netL35 -2.3940722620512824e-13
Rbbr35 netL35 node_2 610.2551678952375
Cbr35 netL35 node_2 -7.430009968873201e-18

* Branch 36
Rabr36 node_1 netRa36 -36.470896460758695
Lbr36 netRa36 netL36 -1.2527753773238529e-13
Rbbr36 netL36 node_2 813.9290073348369
Cbr36 netL36 node_2 -4.357115880614507e-18

* Branch 37
Rabr37 node_1 netRa37 971.4146929189425
Lbr37 netRa37 netL37 9.788608967090214e-13
Rbbr37 netL37 node_2 -4090.0352535072348
Cbr37 netL37 node_2 2.4841024306014845e-19

* Branch 38
Rabr38 node_1 netRa38 -1296.9643370518668
Lbr38 netRa38 netL38 6.960059526687515e-13
Rbbr38 netL38 node_2 2240.4451459359398
Cbr38 netL38 node_2 2.3849347107818596e-19

* Branch 39
Rabr39 node_1 netRa39 -88.31075422567413
Lbr39 netRa39 netL39 -2.060210927051296e-13
Rbbr39 netL39 node_2 563.3857163316061
Cbr39 netL39 node_2 -4.199850883303865e-18

* Branch 40
Rabr40 node_1 netRa40 -51.6785255457787
Lbr40 netRa40 netL40 -1.458824672080668e-13
Rbbr40 netL40 node_2 627.669809837246
Cbr40 netL40 node_2 -4.572060296664842e-18

* Branch 41
Rabr41 node_1 netRa41 8644.436671738453
Lbr41 netRa41 netL41 -2.0187930764058717e-12
Rbbr41 netL41 node_2 -10040.168296132246
Cbr41 netL41 node_2 -2.324523510615043e-20

* Branch 42
Rabr42 node_1 netRa42 132.50765689689158
Lbr42 netRa42 netL42 2.435020651842608e-12
Rbbr42 netL42 node_2 -77633.55144951896
Cbr42 netL42 node_2 2.4544730017904814e-19

* Branch 43
Rabr43 node_1 netRa43 -1563.8531518991506
Lbr43 netRa43 netL43 1.4808282604147074e-12
Rbbr43 netL43 node_2 3712.065606337641
Cbr43 netL43 node_2 2.546428300102819e-19

* Branch 44
Rabr44 node_1 netRa44 11348.749428773379
Lbr44 netRa44 netL44 8.108258120525591e-12
Rbbr44 netL44 node_2 -21857.872479963553
Cbr44 netL44 node_2 3.27202899867656e-20

* Branch 45
Rabr45 node_1 netRa45 -638.8184485192609
Lbr45 netRa45 netL45 5.566847885411315e-13
Rbbr45 netL45 node_2 1842.6115091250708
Cbr45 netL45 node_2 4.723460373170252e-19

* Branch 46
Rabr46 node_1 netRa46 -215.54119563413838
Lbr46 netRa46 netL46 4.97757274242964e-13
Rbbr46 netL46 node_2 3007.2186118907207
Cbr46 netL46 node_2 7.660272209960185e-19

* Branch 47
Rabr47 node_1 netRa47 21568.801887295358
Lbr47 netRa47 netL47 1.075384199777277e-11
Rbbr47 netL47 node_2 -32083.02523463189
Cbr47 netL47 node_2 1.5548257770916648e-20

* Branch 48
Rabr48 node_1 netRa48 372204.7252058415
Lbr48 netRa48 netL48 -3.0980358853001274e-11
Rbbr48 netL48 node_2 -376631.8513707993
Cbr48 netL48 node_2 -2.2098008023464918e-22

* Branch 49
Rabr49 node_1 netRa49 187467.80751448643
Lbr49 netRa49 netL49 1.3471397329167405e-11
Rbbr49 netL49 node_2 -189268.40690595732
Cbr49 netL49 node_2 3.796961100466016e-22

* Branch 50
Rabr50 node_1 netRa50 903458.258688701
Lbr50 netRa50 netL50 5.154000546769364e-11
Rbbr50 netL50 node_2 -909672.2632517148
Cbr50 netL50 node_2 6.271473538986171e-23

* Branch 51
Rabr51 node_1 netRa51 13216176.973375091
Lbr51 netRa51 netL51 -8.146549591876895e-11
Rbbr51 netL51 node_2 -13217695.558979325
Cbr51 netL51 node_2 -4.663481612441336e-25

* Branch 52
Rabr52 node_1 netRa52 159670.80986743682
Lbr52 netRa52 netL52 1.9098107967005588e-11
Rbbr52 netL52 node_2 -164263.8153199847
Cbr52 netL52 node_2 7.282114521854144e-22

* Branch 53
Rabr53 node_1 netRa53 -10179.859007534234
Lbr53 netRa53 netL53 5.505355948515786e-12
Rbbr53 netL53 node_2 15433.909827626776
Cbr53 netL53 node_2 3.5030967706656246e-20

* Branch 54
Rabr54 node_1 netRa54 7432.498174528193
Lbr54 netRa54 netL54 -6.299371917020863e-12
Rbbr54 netL54 node_2 -15382.168319411225
Cbr54 netL54 node_2 -5.508356821297833e-20

* Branch 55
Rabr55 node_1 netRa55 4139.171326619987
Lbr55 netRa55 netL55 8.510194325017899e-12
Rbbr55 netL55 node_2 -40246.108069663605
Cbr55 netL55 node_2 5.111512848703181e-20

* Branch 56
Rabr56 node_1 netRa56 -93133.5377538203
Lbr56 netRa56 netL56 -1.6839031096742724e-11
Rbbr56 netL56 node_2 98955.07292425055
Cbr56 netL56 node_2 -1.8272355265589462e-21

* Branch 57
Rabr57 node_1 netRa57 19986.80818709938
Lbr57 netRa57 netL57 -5.6324220940246185e-12
Rbbr57 netL57 node_2 -23424.308448928445
Cbr57 netL57 node_2 -1.2029718464693292e-20

* Branch 58
Rabr58 node_1 netRa58 -835.8770999860203
Lbr58 netRa58 netL58 7.314994687998328e-12
Rbbr58 netL58 node_2 104652.38984179351
Cbr58 netL58 node_2 8.344770167291228e-20

* Branch 59
Rabr59 node_1 netRa59 -68560.8637613778
Lbr59 netRa59 netL59 2.4910664061260447e-11
Rbbr59 netL59 node_2 82863.31424948243
Cbr59 netL59 node_2 4.3844610318973224e-21

* Branch 60
Rabr60 node_1 netRa60 5261.286365515147
Lbr60 netRa60 netL60 5.277001561525046e-12
Rbbr60 netL60 node_2 -12687.020900022895
Cbr60 netL60 node_2 7.906900832884099e-20

* Branch 61
Rabr61 node_1 netRa61 41036.404616412496
Lbr61 netRa61 netL61 6.618581586347463e-12
Rbbr61 netL61 node_2 -43404.32035041154
Cbr61 netL61 node_2 3.7159253900962146e-21

* Branch 62
Rabr62 node_1 netRa62 -386.5395476194343
Lbr62 netRa62 netL62 -4.358133340616506e-12
Rbbr62 netL62 node_2 23232.200359281516
Cbr62 netL62 node_2 -4.853831424523869e-19

* Branch 63
Rabr63 node_1 netRa63 48949.341431215544
Lbr63 netRa63 netL63 -1.851148207107575e-11
Rbbr63 netL63 node_2 -57616.096483053436
Cbr63 netL63 node_2 -6.5637160786974104e-21

* Branch 64
Rabr64 node_1 netRa64 -481.4123240141128
Lbr64 netRa64 netL64 -4.843529153669744e-12
Rbbr64 netL64 node_2 20811.987285703053
Cbr64 netL64 node_2 -4.834438054024574e-19

* Branch 65
Rabr65 node_1 netRa65 -509.49424784466004
Lbr65 netRa65 netL65 -4.731867442773119e-12
Rbbr65 netL65 node_2 19876.4700948121
Cbr65 netL65 node_2 -4.6726175636526e-19

* Branch 66
Rabr66 node_1 netRa66 20255.21155414322
Lbr66 netRa66 netL66 7.675865661187641e-12
Rbbr66 netL66 node_2 -27183.786955569678
Cbr66 netL66 node_2 1.3940577837544292e-20

* Branch 67
Rabr67 node_1 netRa67 7959.026049510137
Lbr67 netRa67 netL67 5.294846436400066e-12
Rbbr67 netL67 node_2 -15967.36705808941
Cbr67 netL67 node_2 4.166415168774403e-20

* Branch 68
Rabr68 node_1 netRa68 -134.1448438421118
Lbr68 netRa68 netL68 -3.56008572006523e-12
Rbbr68 netL68 node_2 46413.328064614616
Cbr68 netL68 node_2 -5.719351459681622e-19

* Branch 69
Rabr69 node_1 netRa69 9115.634902724565
Lbr69 netRa69 netL69 -1.2569452560400302e-11
Rbbr69 netL69 node_2 -28546.10947029544
Cbr69 netL69 node_2 -4.830296177012301e-20

* Branch 70
Rabr70 node_1 netRa70 389.933518890466
Lbr70 netRa70 netL70 -6.149987389711617e-12
Rbbr70 netL70 node_2 -52857.01662744935
Cbr70 netL70 node_2 -2.9823789701070576e-19

* Branch 71
Rabr71 node_1 netRa71 -56.98291301118493
Lbr71 netRa71 netL71 -5.238052619144044e-12
Rbbr71 netL71 node_2 190562.10981045617
Cbr71 netL71 node_2 -4.838612137460114e-19

* Branch 72
Rabr72 node_1 netRa72 139.31858387276336
Lbr72 netRa72 netL72 -4.795260631392044e-12
Rbbr72 netL72 node_2 -93727.12471269838
Cbr72 netL72 node_2 -3.666184229625398e-19

* Branch 73
Rabr73 node_1 netRa73 10057.296998151698
Lbr73 netRa73 netL73 -1.0707307887775561e-11
Rbbr73 netL73 node_2 -18869.700361922274
Cbr73 netL73 node_2 -5.641717971555052e-20

* Branch 74
Rabr74 node_1 netRa74 2031.4276935512796
Lbr74 netRa74 netL74 -6.427090044106562e-12
Rbbr74 netL74 node_2 -25606.200096379252
Cbr74 netL74 node_2 -1.2353799202878906e-19

* Branch 75
Rabr75 node_1 netRa75 159345.89390248
Lbr75 netRa75 netL75 -5.4145716230732374e-11
Rbbr75 netL75 node_2 -185952.75223546047
Cbr75 netL75 node_2 -1.8273147903632214e-21

* Branch 76
Rabr76 node_1 netRa76 106223.94745995656
Lbr76 netRa76 netL76 2.3641635880036677e-11
Rbbr76 netL76 node_2 -111923.80106235441
Cbr76 netL76 node_2 1.98855524009319e-21

* Branch 77
Rabr77 node_1 netRa77 2218.5007881308093
Lbr77 netRa77 netL77 -4.548834861060225e-12
Rbbr77 netL77 node_2 -8299.747008173075
Cbr77 netL77 node_2 -2.469994749969837e-19

* Branch 78
Rabr78 node_1 netRa78 4291.206550788389
Lbr78 netRa78 netL78 -7.437774224190404e-12
Rbbr78 netL78 node_2 -14668.062658482324
Cbr78 netL78 node_2 -1.1814682751654445e-19

* Branch 79
Rabr79 node_1 netRa79 1998.2619039218323
Lbr79 netRa79 netL79 -3.655808734877788e-12
Rbbr79 netL79 node_2 -6555.282256384778
Cbr79 netL79 node_2 -2.7903819054658453e-19

* Branch 80
Rabr80 node_1 netRa80 531.1660543354797
Lbr80 netRa80 netL80 -3.6953210731448894e-12
Rbbr80 netL80 node_2 -15826.915840509531
Cbr80 netL80 node_2 -4.392603676525071e-19

* Branch 81
Rabr81 node_1 netRa81 3443.09240310078
Lbr81 netRa81 netL81 -5.581721251739968e-12
Rbbr81 netL81 node_2 -11939.601766108113
Cbr81 netL81 node_2 -1.3575548304973188e-19

* Branch 82
Rabr82 node_1 netRa82 19321.20946485749
Lbr82 netRa82 netL82 -8.726854895158264e-12
Rbbr82 netL82 node_2 -21351.03842869138
Cbr82 netL82 node_2 -2.1153337604022513e-20

* Branch 83
Rabr83 node_1 netRa83 2334782.0467978
Lbr83 netRa83 netL83 -1.0790987908347557e-10
Rbbr83 netL83 node_2 -2338481.737378646
Cbr83 netL83 node_2 -1.9764147257327844e-23

* Branch 84
Rabr84 node_1 netRa84 5081.553314168997
Lbr84 netRa84 netL84 -6.678490223015155e-12
Rbbr84 netL84 node_2 -16301.33311958588
Cbr84 netL84 node_2 -8.060726974050976e-20

* Branch 85
Rabr85 node_1 netRa85 16353.690660143346
Lbr85 netRa85 netL85 -9.201706166989245e-12
Rbbr85 netL85 node_2 -21036.84813043193
Cbr85 netL85 node_2 -2.674457373750831e-20

* Branch 86
Rabr86 node_1 netRa86 3362.6224177135555
Lbr86 netRa86 netL86 -3.2263221675966337e-12
Rbbr86 netL86 node_2 -7072.236979921816
Cbr86 netL86 node_2 -1.3564650162923312e-19

* Branch 87
Rabr87 node_1 netRa87 10005.374097753825
Lbr87 netRa87 netL87 -5.630763999587807e-12
Rbbr87 netL87 node_2 -12259.33352888711
Cbr87 netL87 node_2 -4.5900765812624294e-20

* Branch 88
Rabr88 node_1 netRa88 20974.51480091502
Lbr88 netRa88 netL88 -1.1907110195550398e-11
Rbbr88 netL88 node_2 -27801.215703297312
Cbr88 netL88 node_2 -2.041740412674898e-20

* Branch 89
Rabr89 node_1 netRa89 2607.2936333883868
Lbr89 netRa89 netL89 -3.572978566281261e-12
Rbbr89 netL89 node_2 -5659.17644254158
Cbr89 netL89 node_2 -2.4208258495599604e-19

* Branch 90
Rabr90 node_1 netRa90 6568.284298751095
Lbr90 netRa90 netL90 -5.32638349042641e-12
Rbbr90 netL90 node_2 -10329.088223594035
Cbr90 netL90 node_2 -7.849454855364237e-20

* Branch 91
Rabr91 node_1 netRa91 5536.7223898566335
Lbr91 netRa91 netL91 -4.629785113589308e-12
Rbbr91 netL91 node_2 -9587.501936886281
Cbr91 netL91 node_2 -8.719957026539631e-20

* Branch 92
Rabr92 node_1 netRa92 6430.818980063093
Lbr92 netRa92 netL92 -6.64687289035699e-12
Rbbr92 netL92 node_2 -12184.232758976823
Cbr92 netL92 node_2 -8.480759521773152e-20

* Branch 93
Rabr93 node_1 netRa93 389089.12539570755
Lbr93 netRa93 netL93 2.5981464495654496e-11
Rbbr93 netL93 node_2 -391377.7848081184
Cbr93 netL93 node_2 1.7061885999542992e-22

* Branch 94
Rabr94 node_1 netRa94 13221.921850392448
Lbr94 netRa94 netL94 -6.018206939807534e-12
Rbbr94 netL94 node_2 -16950.104868784983
Cbr94 netL94 node_2 -2.684974300261392e-20

* Branch 95
Rabr95 node_1 netRa95 -6609.891706698318
Lbr95 netRa95 netL95 6.416248046142624e-12
Rbbr95 netL95 node_2 21104.829585523064
Cbr95 netL95 node_2 4.5976327172817274e-20

* Branch 96
Rabr96 node_1 netRa96 806633.478788508
Lbr96 netRa96 netL96 2.983366375858232e-11
Rbbr96 netL96 node_2 -807708.4487404717
Cbr96 netL96 node_2 4.5791274293066354e-23

* Branch 97
Rabr97 node_1 netRa97 5488.488092276215
Lbr97 netRa97 netL97 1.3782526147779916e-12
Rbbr97 netL97 node_2 -6552.324993952241
Cbr97 netL97 node_2 3.833437376537022e-20

* Branch 98
Rabr98 node_1 netRa98 227.3026795516643
Lbr98 netRa98 netL98 -1.1433565370580921e-13
Rbbr98 netL98 node_2 -417.6964225306775
Cbr98 netL98 node_2 -1.1836373629096031e-18

* Branch 99
Rabr99 node_1 netRa99 -190.08731344128745
Lbr99 netRa99 netL99 2.5828850384277805e-13
Rbbr99 netL99 node_2 1118.1256337873488
Cbr99 netL99 node_2 1.128903087840525e-18

.ends


* Y'13
.subckt yp13 node_1 node_3
* Branch 0
Rabr0 node_1 netRa0 399.93805556672675
Lbr0 netRa0 netL0 1.651910277578893e-13
Rbbr0 netL0 node_3 -646.9173552745956
Cbr0 netL0 node_3 6.584737557496903e-19

* Branch 1
Rabr1 node_1 netRa1 4476.18768894414
Lbr1 netRa1 netL1 4.865514001834885e-13
Rbbr1 netL1 node_3 -4663.445293900738
Cbr1 netL1 node_3 2.348171186795712e-20

* Branch 2
Rabr2 node_1 netRa2 8116.198793676412
Lbr2 netRa2 netL2 -1.2053250099668384e-12
Rbbr2 netL2 node_3 -8737.049415436175
Cbr2 netL2 node_3 -1.683778695865831e-20

* Branch 3
Rabr3 node_1 netRa3 101.72671211208547
Lbr3 netRa3 netL3 -4.964445135144157e-13
Rbbr3 netL3 node_3 -5406.540752508888
Cbr3 netL3 node_3 -7.170031703710438e-19

* Branch 4
Rabr4 node_1 netRa4 -265.2624396889312
Lbr4 netRa4 netL4 8.183193106731208e-14
Rbbr4 netL4 node_3 351.4771461617258
Cbr4 netL4 node_3 8.643295245310063e-19

* Branch 5
Rabr5 node_1 netRa5 -4557.737175817021
Lbr5 netRa5 netL5 1.3933605631687133e-12
Rbbr5 netL5 node_3 5488.297288462349
Cbr5 netL5 node_3 5.504989752090762e-20

* Branch 6
Rabr6 node_1 netRa6 -17935.2988586583
Lbr6 netRa6 netL6 2.8975221300148818e-12
Rbbr6 netL6 node_3 19424.593978128603
Cbr6 netL6 node_3 8.269906101893293e-21

* Branch 7
Rabr7 node_1 netRa7 -10114.00765606257
Lbr7 netRa7 netL7 2.210898823066605e-12
Rbbr7 netL7 node_3 11191.094430768466
Cbr7 netL7 node_3 1.940039667511203e-20

* Branch 8
Rabr8 node_1 netRa8 -1125.5901013702874
Lbr8 netRa8 netL8 -3.1246138077321283e-13
Rbbr8 netL8 node_3 1418.626462319505
Cbr8 netL8 node_3 -1.9736084455907355e-19

* Branch 9
Rabr9 node_1 netRa9 757.7651931964746
Lbr9 netRa9 netL9 -5.997217582132439e-13
Rbbr9 netL9 node_3 -2040.8486082557993
Cbr9 netL9 node_3 -3.787083967397603e-19

* Branch 10
Rabr10 node_1 netRa10 -15226.065825518524
Lbr10 netRa10 netL10 2.937260745120531e-12
Rbbr10 netL10 node_3 16845.317458883215
Cbr10 netL10 node_3 1.1394340610453182e-20

* Branch 11
Rabr11 node_1 netRa11 -2442.6505099968444
Lbr11 netRa11 netL11 6.912962726161525e-13
Rbbr11 netL11 node_3 3003.835208490254
Cbr11 netL11 node_3 9.352861045034893e-20

* Branch 12
Rabr12 node_1 netRa12 -527.6233822170346
Lbr12 netRa12 netL12 5.753657354994443e-13
Rbbr12 netL12 node_3 1699.4214467461254
Cbr12 netL12 node_3 6.28255859214274e-19

* Branch 13
Rabr13 node_1 netRa13 -102216.70218778489
Lbr13 netRa13 netL13 -4.55099304375019e-12
Rbbr13 netL13 node_3 102785.99384759627
Cbr13 netL13 node_3 -4.335371880419714e-22

* Branch 14
Rabr14 node_1 netRa14 -317.3030695072644
Lbr14 netRa14 netL14 5.356952697688997e-13
Rbbr14 netL14 node_3 1868.7146991324328
Cbr14 netL14 node_3 8.75139071243639e-19

* Branch 15
Rabr15 node_1 netRa15 -262.2162585132483
Lbr15 netRa15 netL15 5.357079082555138e-13
Rbbr15 netL15 node_3 2069.4976385558
Cbr15 netL15 node_3 9.512165468963426e-19

* Branch 16
Rabr16 node_1 netRa16 300088.18615134456
Lbr16 netRa16 netL16 1.027038137958625e-11
Rbbr16 netL16 node_3 -301258.6771791543
Cbr16 netL16 node_3 1.1367597189054373e-22

* Branch 17
Rabr17 node_1 netRa17 -202.8643016326656
Lbr17 netRa17 netL17 5.838569737837363e-13
Rbbr17 netL17 node_3 1907.2514692182717
Cbr17 netL17 node_3 1.4388958221882368e-18

* Branch 18
Rabr18 node_1 netRa18 -61.9602059923413
Lbr18 netRa18 netL18 2.9806921502536526e-13
Rbbr18 netL18 node_3 3892.5042787174543
Cbr18 netL18 node_3 1.1435821496046686e-18

* Branch 19
Rabr19 node_1 netRa19 -32.97699877385237
Lbr19 netRa19 netL19 6.263593019069762e-13
Rbbr19 netL19 node_3 7888.235196079105
Cbr19 netL19 node_3 1.8793197516850748e-18

* Branch 20
Rabr20 node_1 netRa20 -168.89921608745846
Lbr20 netRa20 netL20 5.573514930315672e-13
Rbbr20 netL20 node_3 2663.119269669761
Cbr20 netL20 node_3 1.18186274839003e-18

* Branch 21
Rabr21 node_1 netRa21 -74.03180630113316
Lbr21 netRa21 netL21 5.863791626617302e-13
Rbbr21 netL21 node_3 4006.9167719188586
Cbr21 netL21 node_3 1.7806259976772892e-18

* Branch 22
Rabr22 node_1 netRa22 -202911740.5805401
Lbr22 netRa22 netL22 -2.2546556583098137e-10
Rbbr22 netL22 node_3 202912353.8869405
Cbr22 netL22 node_3 -5.4760986685630744e-27

* Branch 23
Rabr23 node_1 netRa23 182.07441937642162
Lbr23 netRa23 netL23 8.483877997323419e-13
Rbbr23 netL23 node_3 -2831.4878508603133
Cbr23 netL23 node_3 1.7592734391879437e-18

* Branch 24
Rabr24 node_1 netRa24 -12.391793550861086
Lbr24 netRa24 netL24 6.788439883149488e-13
Rbbr24 netL24 node_3 16734.26117297341
Cbr24 netL24 node_3 1.904946922437278e-18

* Branch 25
Rabr25 node_1 netRa25 -6961.874758298142
Lbr25 netRa25 netL25 2.8822637014961855e-12
Rbbr25 netL25 node_3 10657.51269300898
Cbr25 netL25 node_3 3.8644857102647934e-20

* Branch 26
Rabr26 node_1 netRa26 -128.05883175882468
Lbr26 netRa26 netL26 5.689848609862655e-13
Rbbr26 netL26 node_3 2573.9625950970594
Cbr26 netL26 node_3 1.6387737895841431e-18

* Branch 27
Rabr27 node_1 netRa27 -122.0922912623511
Lbr27 netRa27 netL27 1.0510648705554973e-12
Rbbr27 netL27 node_3 4452.48113261231
Cbr27 netL27 node_3 1.7529983879338707e-18

* Branch 28
Rabr28 node_1 netRa28 38789.349482970654
Lbr28 netRa28 netL28 4.888867655923921e-12
Rbbr28 netL28 node_3 -40191.59135135048
Cbr28 netL28 node_3 3.140298477583059e-21

* Branch 29
Rabr29 node_1 netRa29 -191.45954264361873
Lbr29 netRa29 netL29 5.495053613615792e-13
Rbbr29 netL29 node_3 2656.605069350042
Cbr29 netL29 node_3 1.0471656261035982e-18

* Branch 30
Rabr30 node_1 netRa30 -141.20605319630494
Lbr30 netRa30 netL30 5.594778807385958e-13
Rbbr30 netL30 node_3 3110.678098629599
Cbr30 netL30 node_3 1.220532141249798e-18

* Branch 31
Rabr31 node_1 netRa31 -425.34429685482843
Lbr31 netRa31 netL31 -4.3124633475115166e-13
Rbbr31 netL31 node_3 1545.5091186928892
Cbr31 netL31 node_3 -6.626721209398794e-19

* Branch 32
Rabr32 node_1 netRa32 313.7555176595352
Lbr32 netRa32 netL32 9.355189916843174e-13
Rbbr32 netL32 node_3 -2077.90596128577
Cbr32 netL32 node_3 1.4785902070511907e-18

* Branch 33
Rabr33 node_1 netRa33 -578.1369665237935
Lbr33 netRa33 netL33 -8.287821325213738e-13
Rbbr33 netL33 node_3 4710.957816908979
Cbr33 netL33 node_3 -3.081994575274113e-19

* Branch 34
Rabr34 node_1 netRa34 -83.5449552858749
Lbr34 netRa34 netL34 5.764830887959441e-13
Rbbr34 netL34 node_3 4989.39022017772
Cbr34 netL34 node_3 1.3066639908698835e-18

* Branch 35
Rabr35 node_1 netRa35 -1160.5168188258203
Lbr35 netRa35 netL35 6.993741737242146e-13
Rbbr35 netL35 node_3 2034.9046934562077
Cbr35 netL35 node_3 2.9473364276665127e-19

* Branch 36
Rabr36 node_1 netRa36 2.734965693957903
Lbr36 netRa36 netL36 6.777996797519927e-13
Rbbr36 netL36 node_3 153229.93566524473
Cbr36 netL36 node_3 2.1320638767793113e-18

* Branch 37
Rabr37 node_1 netRa37 -718.5836777054363
Lbr37 netRa37 netL37 -1.7863253159477074e-12
Rbbr37 netL37 node_3 3304.1338784448376
Cbr37 netL37 node_3 -7.656221339477291e-19

* Branch 38
Rabr38 node_1 netRa38 497.0875273159017
Lbr38 netRa38 netL38 2.3181584798996216e-12
Rbbr38 netL38 node_3 -34339.015117905765
Cbr38 netL38 node_3 1.4035391328972294e-19

* Branch 39
Rabr39 node_1 netRa39 4066000.956928218
Lbr39 netRa39 netL39 1.6506050732617232e-10
Rbbr39 netL39 node_3 -4073530.3062922894
Cbr39 netL39 node_3 9.968392042491645e-24

* Branch 40
Rabr40 node_1 netRa40 2425.782454355772
Lbr40 netRa40 netL40 1.6004679131063655e-12
Rbbr40 netL40 node_3 -5567.749820211374
Cbr40 netL40 node_3 1.1903257292080075e-19

* Branch 41
Rabr41 node_1 netRa41 107.51174555752745
Lbr41 netRa41 netL41 7.610660130273319e-13
Rbbr41 netL41 node_3 -6958.467110444396
Cbr41 netL41 node_3 1.0683243254429985e-18

* Branch 42
Rabr42 node_1 netRa42 -3857.970050664179
Lbr42 netRa42 netL42 1.0239628374329322e-12
Rbbr42 netL42 node_3 4554.080542597762
Cbr42 netL42 node_3 5.818042947887518e-20

* Branch 43
Rabr43 node_1 netRa43 227.0868229263117
Lbr43 netRa43 netL43 1.380730571438887e-12
Rbbr43 netL43 node_3 -24031.473113056185
Cbr43 netL43 node_3 2.6310670859236517e-19

* Branch 44
Rabr44 node_1 netRa44 80859.04038833955
Lbr44 netRa44 netL44 -1.8418919653987138e-11
Rbbr44 netL44 node_3 -83155.68038304689
Cbr44 netL44 node_3 -2.7356285461352202e-21

* Branch 45
Rabr45 node_1 netRa45 -286.51069743115227
Lbr45 netRa45 netL45 5.496321589326636e-13
Rbbr45 netL45 node_3 808.4376986637295
Cbr45 netL45 node_3 2.346858319512148e-18

* Branch 46
Rabr46 node_1 netRa46 -3354.073549330745
Lbr46 netRa46 netL46 -1.0621883957324274e-11
Rbbr46 netL46 node_3 43265.37313996582
Cbr46 netL46 node_3 -7.454933515990913e-20

* Branch 47
Rabr47 node_1 netRa47 125.00695244771707
Lbr47 netRa47 netL47 -2.6080099302474605e-13
Rbbr47 netL47 node_3 -1674.844535749034
Cbr47 netL47 node_3 -1.2317515719282134e-18

* Branch 48
Rabr48 node_1 netRa48 -1614.9934139046543
Lbr48 netRa48 netL48 -2.5845782378010845e-12
Rbbr48 netL48 node_3 3652.5897003102673
Cbr48 netL48 node_3 -4.399911160751773e-19

* Branch 49
Rabr49 node_1 netRa49 -524.9811420872594
Lbr49 netRa49 netL49 1.505236692345846e-12
Rbbr49 netL49 node_3 3058.985682755071
Cbr49 netL49 node_3 9.30326133852985e-19

* Branch 50
Rabr50 node_1 netRa50 -14218.268601274185
Lbr50 netRa50 netL50 -8.857594059542442e-12
Rbbr50 netL50 node_3 22946.209601984712
Cbr50 netL50 node_3 -2.719162014568248e-20

* Branch 51
Rabr51 node_1 netRa51 -3517.690575783094
Lbr51 netRa51 netL51 -3.3629663855193193e-12
Rbbr51 netL51 node_3 7386.649469947278
Cbr51 netL51 node_3 -1.2973111009568104e-19

* Branch 52
Rabr52 node_1 netRa52 6354.290147374493
Lbr52 netRa52 netL52 5.420805791592377e-12
Rbbr52 netL52 node_3 -17163.589097844433
Cbr52 netL52 node_3 4.979774064284513e-20

* Branch 53
Rabr53 node_1 netRa53 -3211.3166148633786
Lbr53 netRa53 netL53 2.7811798811598294e-12
Rbbr53 netL53 node_3 9493.421843937791
Cbr53 netL53 node_3 9.106038002302316e-20

* Branch 54
Rabr54 node_1 netRa54 -519.1704032540396
Lbr54 netRa54 netL54 4.145648815302462e-12
Rbbr54 netL54 node_3 87534.08575833886
Cbr54 netL54 node_3 8.985206547728025e-20

* Branch 55
Rabr55 node_1 netRa55 -22413.786054228727
Lbr55 netRa55 netL55 -1.793256208970298e-11
Rbbr55 netL55 node_3 28758.749064332966
Cbr55 netL55 node_3 -2.7857961344376257e-20

* Branch 56
Rabr56 node_1 netRa56 -9848.43677553974
Lbr56 netRa56 netL56 -1.1623845486189636e-11
Rbbr56 netL56 node_3 16249.52545461652
Cbr56 netL56 node_3 -7.275583660297246e-20

* Branch 57
Rabr57 node_1 netRa57 -13455.314832242198
Lbr57 netRa57 netL57 -1.2679887062351811e-11
Rbbr57 netL57 node_3 28764.41106802511
Cbr57 netL57 node_3 -3.279623503081049e-20

* Branch 58
Rabr58 node_1 netRa58 -1060340.127491106
Lbr58 netRa58 netL58 1.6582593008553795e-10
Rbbr58 netL58 node_3 1071170.7993329733
Cbr58 netL58 node_3 1.4597568014434174e-22

* Branch 59
Rabr59 node_1 netRa59 -74345.67789052027
Lbr59 netRa59 netL59 -8.695681403500898e-11
Rbbr59 netL59 node_3 230601.57825136048
Cbr59 netL59 node_3 -5.0776303527446165e-21

* Branch 60
Rabr60 node_1 netRa60 378937.7484031683
Lbr60 netRa60 netL60 -2.0552419574205954e-10
Rbbr60 netL60 node_3 -458287.9039330575
Cbr60 netL60 node_3 -1.1829216056322199e-21

* Branch 61
Rabr61 node_1 netRa61 12230.150965646653
Lbr61 netRa61 netL61 -1.7613318806386517e-11
Rbbr61 netL61 node_3 -39678.50968158748
Cbr61 netL61 node_3 -3.6259338184429513e-20

* Branch 62
Rabr62 node_1 netRa62 -2722236.1995962705
Lbr62 netRa62 netL62 3.149499833222646e-10
Rbbr62 netL62 node_3 2749292.5010153963
Cbr62 netL62 node_3 4.207873804292648e-23

* Branch 63
Rabr63 node_1 netRa63 -16701.1357672465
Lbr63 netRa63 netL63 -2.478502240889619e-11
Rbbr63 netL63 node_3 45180.59845567062
Cbr63 netL63 node_3 -3.2872495213698535e-20

* Branch 64
Rabr64 node_1 netRa64 -91465.17238872804
Lbr64 netRa64 netL64 8.373491078151097e-11
Rbbr64 netL64 node_3 153194.44283036297
Cbr64 netL64 node_3 5.973499650536987e-21

* Branch 65
Rabr65 node_1 netRa65 357686.4032854409
Lbr65 netRa65 netL65 9.13642071885978e-11
Rbbr65 netL65 node_3 -391459.38714078505
Cbr65 netL65 node_3 6.52576215547816e-22

* Branch 66
Rabr66 node_1 netRa66 -9034.767922946094
Lbr66 netRa66 netL66 2.885478847735536e-11
Rbbr66 netL66 node_3 45365.752103987164
Cbr66 netL66 node_3 7.032398191973406e-20

* Branch 67
Rabr67 node_1 netRa67 249797.45858933005
Lbr67 netRa67 netL67 2.3015375006996674e-10
Rbbr67 netL67 node_3 -565911.7724955818
Cbr67 netL67 node_3 1.6285984121284844e-21

* Branch 68
Rabr68 node_1 netRa68 -440134.5153571677
Lbr68 netRa68 netL68 1.1609370688744101e-10
Rbbr68 netL68 node_3 465794.83959805116
Cbr68 netL68 node_3 5.66229698901179e-22

* Branch 69
Rabr69 node_1 netRa69 14706826.126101395
Lbr69 netRa69 netL69 5.246567871583091e-10
Rbbr69 netL69 node_3 -14737243.084582895
Cbr69 netL69 node_3 2.420722128311739e-24

* Branch 70
Rabr70 node_1 netRa70 -30647.80307678151
Lbr70 netRa70 netL70 -3.484715904460165e-11
Rbbr70 netL70 node_3 112395.75917038362
Cbr70 netL70 node_3 -1.0119769736082296e-20

* Branch 71
Rabr71 node_1 netRa71 -13515.47958249684
Lbr71 netRa71 netL71 -3.239668507414866e-11
Rbbr71 netL71 node_3 62004.502988120934
Cbr71 netL71 node_3 -3.868646921229621e-20

* Branch 72
Rabr72 node_1 netRa72 75498.03028299888
Lbr72 netRa72 netL72 -5.192987570384009e-11
Rbbr72 netL72 node_3 -143738.2762885616
Cbr72 netL72 node_3 -4.7843710334423676e-21

* Branch 73
Rabr73 node_1 netRa73 -12731.75255474266
Lbr73 netRa73 netL73 8.559186293907941e-11
Rbbr73 netL73 node_3 513084.97747974994
Cbr73 netL73 node_3 1.3077811864468265e-20

* Branch 74
Rabr74 node_1 netRa74 -29241.66707089115
Lbr74 netRa74 netL74 4.94365555197482e-11
Rbbr74 netL74 node_3 104867.90847279219
Cbr74 netL74 node_3 1.61174357355722e-20

* Branch 75
Rabr75 node_1 netRa75 11035.741779748052
Lbr75 netRa75 netL75 5.390717254578808e-11
Rbbr75 netL75 node_3 -451175.7236563157
Cbr75 netL75 node_3 1.0833596957381712e-20

* Branch 76
Rabr76 node_1 netRa76 -135512.83386851035
Lbr76 netRa76 netL76 -7.402614285941694e-11
Rbbr76 netL76 node_3 206868.19745334884
Cbr76 netL76 node_3 -2.640715968772765e-21

* Branch 77
Rabr77 node_1 netRa77 257463.69705420523
Lbr77 netRa77 netL77 -1.194376674344107e-10
Rbbr77 netL77 node_3 -357879.5070555878
Cbr77 netL77 node_3 -1.2962252655980252e-21

* Branch 78
Rabr78 node_1 netRa78 -1754.8376047607067
Lbr78 netRa78 netL78 -7.435745639916701e-11
Rbbr78 netL78 node_3 2154148.2726473175
Cbr78 netL78 node_3 -1.9701874158189738e-20

* Branch 79
Rabr79 node_1 netRa79 -5388.082042079682
Lbr79 netRa79 netL79 7.701439694567752e-11
Rbbr79 netL79 node_3 723483.6614024995
Cbr79 netL79 node_3 1.975322604292801e-20

* Branch 80
Rabr80 node_1 netRa80 24736.661798549205
Lbr80 netRa80 netL80 -4.5423599000735473e-11
Rbbr80 netL80 node_3 -128132.5943962454
Cbr80 netL80 node_3 -1.4331117915418528e-20

* Branch 81
Rabr81 node_1 netRa81 -87007.09266323024
Lbr81 netRa81 netL81 4.937188721705374e-11
Rbbr81 netL81 node_3 113326.89893733885
Cbr81 netL81 node_3 5.007127541567701e-21

* Branch 82
Rabr82 node_1 netRa82 -8063108.28807664
Lbr82 netRa82 netL82 5.38129274597605e-10
Rbbr82 netL82 node_3 8124776.911928087
Cbr82 netL82 node_3 8.214330399677914e-24

* Branch 83
Rabr83 node_1 netRa83 -1037870.9563077653
Lbr83 netRa83 netL83 -2.352329699158334e-10
Rbbr83 netL83 node_3 1112715.822814586
Cbr83 netL83 node_3 -2.0369137643439929e-22

* Branch 84
Rabr84 node_1 netRa84 -1653002.9079265124
Lbr84 netRa84 netL84 2.3883740463088683e-10
Rbbr84 netL84 node_3 1689120.3250563235
Cbr84 netL84 node_3 8.553940775354375e-23

* Branch 85
Rabr85 node_1 netRa85 -1711670.9549001171
Lbr85 netRa85 netL85 4.6110025455685095e-10
Rbbr85 netL85 node_3 1942860.3053938253
Cbr85 netL85 node_3 1.3865104538392648e-22

* Branch 86
Rabr86 node_1 netRa86 7280499048.461896
Lbr86 netRa86 netL86 1.3641501770012138e-08
Rbbr86 netL86 node_3 -7280532805.0780115
Cbr86 netL86 node_3 2.5735817597207515e-28

* Branch 87
Rabr87 node_1 netRa87 81315.84502179541
Lbr87 netRa87 netL87 -4.49944908889338e-11
Rbbr87 netL87 node_3 -143434.81272305807
Cbr87 netL87 node_3 -3.8573915017035e-21

* Branch 88
Rabr88 node_1 netRa88 -683687.0117867832
Lbr88 netRa88 netL88 2.949028853185057e-10
Rbbr88 netL88 node_3 939486.9375639132
Cbr88 netL88 node_3 4.590943822190674e-22

* Branch 89
Rabr89 node_1 netRa89 -17947.172352426274
Lbr89 netRa89 netL89 3.050067122168343e-11
Rbbr89 netL89 node_3 68450.78768803916
Cbr89 netL89 node_3 2.4820909285831626e-20

* Branch 90
Rabr90 node_1 netRa90 359394.7584853014
Lbr90 netRa90 netL90 1.6795297686413078e-10
Rbbr90 netL90 node_3 -513264.04285211564
Cbr90 netL90 node_3 9.105733109716915e-22

* Branch 91
Rabr91 node_1 netRa91 -140302.91712423798
Lbr91 netRa91 netL91 4.511719092890651e-11
Rbbr91 netL91 node_3 154960.61705220488
Cbr91 netL91 node_3 2.07502880805208e-21

* Branch 92
Rabr92 node_1 netRa92 9344.698105590853
Lbr92 netRa92 netL92 1.510935751666023e-11
Rbbr92 netL92 node_3 -62286.34457568919
Cbr92 netL92 node_3 2.5969437611941735e-20

* Branch 93
Rabr93 node_1 netRa93 611985.5953015708
Lbr93 netRa93 netL93 7.647992896475671e-11
Rbbr93 netL93 node_3 -632186.7460497809
Cbr93 netL93 node_3 1.9768549121177467e-22

* Branch 94
Rabr94 node_1 netRa94 -10744.627671151973
Lbr94 netRa94 netL94 -1.6150720687846678e-11
Rbbr94 netL94 node_3 43823.22548665498
Cbr94 netL94 node_3 -3.4317847666879746e-20

* Branch 95
Rabr95 node_1 netRa95 23346.620243439756
Lbr95 netRa95 netL95 -2.0117943966881866e-11
Rbbr95 netL95 node_3 -65609.20621479608
Cbr95 netL95 node_3 -1.3127216360242349e-20

* Branch 96
Rabr96 node_1 netRa96 65873.94332416392
Lbr96 netRa96 netL96 -2.7258366764215506e-11
Rbbr96 netL96 node_3 -92766.82390787534
Cbr96 netL96 node_3 -4.4594403923239635e-21

* Branch 97
Rabr97 node_1 netRa97 94945.46234044811
Lbr97 netRa97 netL97 -4.11296533444881e-11
Rbbr97 netL97 node_3 -134457.65695778705
Cbr97 netL97 node_3 -3.220711897941488e-21

* Branch 98
Rabr98 node_1 netRa98 -110.11933558740924
Lbr98 netRa98 netL98 6.163024806447084e-13
Rbbr98 netL98 node_3 9183.069681130513
Cbr98 netL98 node_3 5.5750636595264305e-19

* Branch 99
Rabr99 node_1 netRa99 123080.37708135683
Lbr99 netRa99 netL99 -2.9446710226876348e-12
Rbbr99 netL99 node_3 -123327.23714292314
Cbr99 netL99 node_3 -1.936912559939517e-22

.ends


* Y'14
.subckt yp14 node_1 node_4
* Branch 0
Rabr0 node_1 netRa0 -644.8228390438431
Lbr0 netRa0 netL0 2.1398670101037786e-13
Rbbr0 netL0 node_4 883.431971930877
Cbr0 netL0 node_4 3.655607026802236e-19

* Branch 1
Rabr1 node_1 netRa1 912.98410381908
Lbr1 netRa1 netL1 2.2664133225208223e-13
Rbbr1 netL1 node_4 -1111.0822836677164
Cbr1 netL1 node_4 2.2791213216641855e-19

* Branch 2
Rabr2 node_1 netRa2 378.458165809748
Lbr2 netRa2 netL2 -6.667918550102573e-14
Rbbr2 netL2 node_4 -418.46660490768915
Cbr2 netL2 node_4 -4.1577430779990005e-19

* Branch 3
Rabr3 node_1 netRa3 -28.670908096235678
Lbr3 netRa3 netL3 2.632073993288762e-14
Rbbr3 netL3 node_4 93.38579841360728
Cbr3 netL3 node_4 9.250872622247668e-18

* Branch 4
Rabr4 node_1 netRa4 -14.636712535005504
Lbr4 netRa4 netL4 2.431189435077642e-14
Rbbr4 netL4 node_4 118.6440258376462
Cbr4 netL4 node_4 1.2670614676405491e-17

* Branch 5
Rabr5 node_1 netRa5 -49.88377514692712
Lbr5 netRa5 netL5 3.5004020465414787e-14
Rbbr5 netL5 node_4 129.8682602409046
Cbr5 netL5 node_4 5.186458352796558e-18

* Branch 6
Rabr6 node_1 netRa6 -0.17111764214529498
Lbr6 netRa6 netL6 2.313201277377136e-14
Rbbr6 netL6 node_4 1016.0504105233654
Cbr6 netL6 node_4 1.5195734987150867e-17

* Branch 7
Rabr7 node_1 netRa7 -49.720463185913424
Lbr7 netRa7 netL7 -2.9720570386241007e-14
Rbbr7 netL7 node_4 100.58974765787714
Cbr7 netL7 node_4 -6.126140165206444e-18

* Branch 8
Rabr8 node_1 netRa8 18088.284455805937
Lbr8 netRa8 netL8 -6.401470266125119e-13
Rbbr8 netL8 node_4 -18152.13692506125
Cbr8 netL8 node_4 -1.94639470169859e-21

* Branch 9
Rabr9 node_1 netRa9 -34.52430970770706
Lbr9 netRa9 netL9 -1.9558860576910455e-14
Rbbr9 netL9 node_4 65.75595465615343
Cbr9 netL9 node_4 -8.794146381333761e-18

* Branch 10
Rabr10 node_1 netRa10 -374.07074386033594
Lbr10 netRa10 netL10 -9.725453926970653e-14
Rbbr10 netL10 node_4 431.30648068701623
Cbr10 netL10 node_4 -6.081665099099981e-19

* Branch 11
Rabr11 node_1 netRa11 -13336.897594380402
Lbr11 netRa11 netL11 1.208716046226364e-12
Rbbr11 netL11 node_4 13607.808147343798
Cbr11 netL11 node_4 6.642186529318227e-21

* Branch 12
Rabr12 node_1 netRa12 -3155.9885585917323
Lbr12 netRa12 netL12 -4.3984848474584714e-13
Rbbr12 netL12 node_4 3307.1121347065723
Cbr12 netL12 node_4 -4.23132244214189e-20

* Branch 13
Rabr13 node_1 netRa13 -1942.8161534478315
Lbr13 netRa13 netL13 -7.040834944332846e-13
Rbbr13 netL13 node_4 2785.04384865697
Cbr13 netL13 node_4 -1.3143625354318318e-19

* Branch 14
Rabr14 node_1 netRa14 2237.538134742306
Lbr14 netRa14 netL14 3.254514592324128e-13
Rbbr14 netL14 node_4 -2379.939153710632
Cbr14 netL14 node_4 6.135639833242439e-20

* Branch 15
Rabr15 node_1 netRa15 18441.619389018117
Lbr15 netRa15 netL15 8.701552889966006e-13
Rbbr15 netL15 node_4 -18561.702330897428
Cbr15 netL15 node_4 2.5451971673666205e-21

* Branch 16
Rabr16 node_1 netRa16 -194.29249821165155
Lbr16 netRa16 netL16 1.3097517418763026e-13
Rbbr16 netL16 node_4 394.019501483195
Cbr16 netL16 node_4 1.6811384614089268e-18

* Branch 17
Rabr17 node_1 netRa17 -97.09114139900433
Lbr17 netRa17 netL17 1.017844419626014e-13
Rbbr17 netL17 node_4 359.51678188644786
Cbr17 netL17 node_4 2.8472499462022763e-18

* Branch 18
Rabr18 node_1 netRa18 -734.1516476740865
Lbr18 netRa18 netL18 -2.3521541557229895e-13
Rbbr18 netL18 node_4 921.2105158813831
Cbr18 netL18 node_4 -3.502384863098941e-19

* Branch 19
Rabr19 node_1 netRa19 -11.958625717934382
Lbr19 netRa19 netL19 -9.775338652355323e-14
Rbbr19 netL19 node_4 1785.0425001703015
Cbr19 netL19 node_4 -5.497367819264466e-18

* Branch 20
Rabr20 node_1 netRa20 201.92915442280074
Lbr20 netRa20 netL20 -2.3571267129530223e-13
Rbbr20 netL20 node_4 -1018.819230224345
Cbr20 netL20 node_4 -1.1198704010545803e-18

* Branch 21
Rabr21 node_1 netRa21 -5.526227931359877
Lbr21 netRa21 netL21 -7.700287691902764e-14
Rbbr21 netL21 node_4 2414.0340938496997
Cbr21 netL21 node_4 -7.46574722870242e-18

* Branch 22
Rabr22 node_1 netRa22 -4.236681938865182
Lbr22 netRa22 netL22 -4.801485990461667e-14
Rbbr22 netL22 node_4 572.9366656541545
Cbr22 netL22 node_4 -2.4192862018004857e-17

* Branch 23
Rabr23 node_1 netRa23 -546.9246211743334
Lbr23 netRa23 netL23 1.714662106828016e-13
Rbbr23 netL23 node_4 661.7470586602029
Cbr23 netL23 node_4 4.714175669395005e-19

* Branch 24
Rabr24 node_1 netRa24 9.0190100188559
Lbr24 netRa24 netL24 -3.856069186166144e-14
Rbbr24 netL24 node_4 -177.16677796047261
Cbr24 netL24 node_4 -2.264083034835337e-17

* Branch 25
Rabr25 node_1 netRa25 -5.133404650062858
Lbr25 netRa25 netL25 -5.202566889214636e-14
Rbbr25 netL25 node_4 483.0365110260438
Cbr25 netL25 node_4 -2.4353259052167422e-17

* Branch 26
Rabr26 node_1 netRa26 -2.6473951558080424
Lbr26 netRa26 netL26 -5.481014136226209e-14
Rbbr26 netL26 node_4 2330.5073422976357
Cbr26 netL26 node_4 -1.2358036782035358e-17

* Branch 27
Rabr27 node_1 netRa27 -1.1763280766955844
Lbr27 netRa27 netL27 -4.633769835839776e-14
Rbbr27 netL27 node_4 3361.0997820757607
Cbr27 netL27 node_4 -2.2908501005351853e-17

* Branch 28
Rabr28 node_1 netRa28 -263.49938435499985
Lbr28 netRa28 netL28 -2.6857676150173573e-13
Rbbr28 netL28 node_4 814.9081349588358
Cbr28 netL28 node_4 -1.2664667394207948e-18

* Branch 29
Rabr29 node_1 netRa29 -39.7603375294024
Lbr29 netRa29 netL29 -7.971590685753722e-14
Rbbr29 netL29 node_4 225.5842679613942
Cbr29 netL29 node_4 -9.097516369349962e-18

* Branch 30
Rabr30 node_1 netRa30 268.8883084311438
Lbr30 netRa30 netL30 -2.480677316775574e-13
Rbbr30 netL30 node_4 -815.0706693072165
Cbr30 netL30 node_4 -1.1201498833987022e-18

* Branch 31
Rabr31 node_1 netRa31 0.8401013331765004
Lbr31 netRa31 netL31 -4.370550925169543e-14
Rbbr31 netL31 node_4 -1482.212410129192
Cbr31 netL31 node_4 -2.2358316781557428e-17

* Branch 32
Rabr32 node_1 netRa32 1785.2626568574315
Lbr32 netRa32 netL32 -9.26743891887414e-13
Rbbr32 netL32 node_4 -3414.185401558983
Cbr32 netL32 node_4 -1.5121554659343788e-19

* Branch 33
Rabr33 node_1 netRa33 13.636205816109428
Lbr33 netRa33 netL33 -5.100925938499105e-14
Rbbr33 netL33 node_4 -111.78810167623307
Cbr33 netL33 node_4 -3.233490316191904e-17

* Branch 34
Rabr34 node_1 netRa34 -4.450161829441548
Lbr34 netRa34 netL34 -7.558944563205361e-14
Rbbr34 netL34 node_4 2526.271254737357
Cbr34 netL34 node_4 -7.954456076344518e-18

* Branch 35
Rabr35 node_1 netRa35 -11.022793544353643
Lbr35 netRa35 netL35 -5.960407481142523e-14
Rbbr35 netL35 node_4 225.89824215756886
Cbr35 netL35 node_4 -2.5162798028004212e-17

* Branch 36
Rabr36 node_1 netRa36 10.586726770007488
Lbr36 netRa36 netL36 -6.318579445480859e-14
Rbbr36 netL36 node_4 -453.65383549594105
Cbr36 netL36 node_4 -1.2493735740409301e-17

* Branch 37
Rabr37 node_1 netRa37 -5.805275937081227
Lbr37 netRa37 netL37 -5.842011129623426e-14
Rbbr37 netL37 node_4 914.7560974466388
Cbr37 netL37 node_4 -1.2058589309687057e-17

* Branch 38
Rabr38 node_1 netRa38 45913.713016128895
Lbr38 netRa38 netL38 -6.4843230590160596e-12
Rbbr38 netL38 node_4 -48766.43412327034
Cbr38 netL38 node_4 -2.892670232764642e-21

* Branch 39
Rabr39 node_1 netRa39 -13.001545874053814
Lbr39 netRa39 netL39 -6.140891942737361e-14
Rbbr39 netL39 node_4 198.99000989810756
Cbr39 netL39 node_4 -2.4645249071780732e-17

* Branch 40
Rabr40 node_1 netRa40 18257.0066919746
Lbr40 netRa40 netL40 -7.175699283537035e-12
Rbbr40 netL40 node_4 -24893.550935108244
Cbr40 netL40 node_4 -1.574438133811996e-20

* Branch 41
Rabr41 node_1 netRa41 -21.85924042079633
Lbr41 netRa41 netL41 -7.500902865027618e-14
Rbbr41 netL41 node_4 167.2702927279277
Cbr41 netL41 node_4 -2.098601477732831e-17

* Branch 42
Rabr42 node_1 netRa42 -1479.8615650495294
Lbr42 netRa42 netL42 -1.1960154524369769e-12
Rbbr42 netL42 node_4 4708.150530596769
Cbr42 netL42 node_4 -1.725464288966709e-19

* Branch 43
Rabr43 node_1 netRa43 -2.5477792511837567
Lbr43 netRa43 netL43 -4.99485792007326e-14
Rbbr43 netL43 node_4 775.5002873103809
Cbr43 netL43 node_4 -2.848367329802999e-17

* Branch 44
Rabr44 node_1 netRa44 -68.749647062703
Lbr44 netRa44 netL44 -1.0827827305142113e-13
Rbbr44 netL44 node_4 270.95464288944305
Cbr44 netL44 node_4 -5.864843844210488e-18

* Branch 45
Rabr45 node_1 netRa45 3846.7163094739753
Lbr45 netRa45 netL45 5.568602770661776e-13
Rbbr45 netL45 node_4 -4064.7216698142233
Cbr45 netL45 node_4 3.56409863275102e-20

* Branch 46
Rabr46 node_1 netRa46 16.226681472899568
Lbr46 netRa46 netL46 -4.2782789039516445e-14
Rbbr46 netL46 node_4 -72.46156820252176
Cbr46 netL46 node_4 -3.5913317547612484e-17

* Branch 47
Rabr47 node_1 netRa47 -236.34186958444673
Lbr47 netRa47 netL47 -4.842757856062195e-13
Rbbr47 netL47 node_4 812.9982169341384
Cbr47 netL47 node_4 -2.54383181212241e-18

* Branch 48
Rabr48 node_1 netRa48 -405.78262805212154
Lbr48 netRa48 netL48 2.2638446216011297e-13
Rbbr48 netL48 node_4 759.6890244985004
Cbr48 netL48 node_4 7.326250101078917e-19

* Branch 49
Rabr49 node_1 netRa49 17861.59758102973
Lbr49 netRa49 netL49 -3.103516081241692e-12
Rbbr49 netL49 node_4 -18182.904667081468
Cbr49 netL49 node_4 -9.550708669821867e-21

* Branch 50
Rabr50 node_1 netRa50 -30.58312460860991
Lbr50 netRa50 netL50 -7.795499793571453e-14
Rbbr50 netL50 node_4 296.7387790313879
Cbr50 netL50 node_4 -8.64014471576844e-18

* Branch 51
Rabr51 node_1 netRa51 -600.074892672273
Lbr51 netRa51 netL51 -5.523451977701148e-13
Rbbr51 netL51 node_4 1213.9900178886478
Cbr51 netL51 node_4 -7.597061119742014e-19

* Branch 52
Rabr52 node_1 netRa52 904.3234943521918
Lbr52 netRa52 netL52 7.406097722478193e-13
Rbbr52 netL52 node_4 -1707.3732448755663
Cbr52 netL52 node_4 4.802329859394199e-19

* Branch 53
Rabr53 node_1 netRa53 1657.8078507276753
Lbr53 netRa53 netL53 5.204813402694056e-13
Rbbr53 netL53 node_4 -2058.97233042227
Cbr53 netL53 node_4 1.5254628959293217e-19

* Branch 54
Rabr54 node_1 netRa54 10.241770674603082
Lbr54 netRa54 netL54 2.0938276448376823e-13
Rbbr54 netL54 node_4 -2155.0811180211485
Cbr54 netL54 node_4 9.6675073420649e-18

* Branch 55
Rabr55 node_1 netRa55 -134.20187110265155
Lbr55 netRa55 netL55 -3.251784715641891e-13
Rbbr55 netL55 node_4 1148.268011892502
Cbr55 netL55 node_4 -2.1147467221585633e-18

* Branch 56
Rabr56 node_1 netRa56 -960.5015385029984
Lbr56 netRa56 netL56 -8.271091446015354e-13
Rbbr56 netL56 node_4 1468.8875943816697
Cbr56 netL56 node_4 -5.866776711591325e-19

* Branch 57
Rabr57 node_1 netRa57 254.325878945563
Lbr57 netRa57 netL57 7.539502550243952e-13
Rbbr57 netL57 node_4 -1245.5470690867887
Cbr57 netL57 node_4 2.386080869805903e-18

* Branch 58
Rabr58 node_1 netRa58 -779.6495548368741
Lbr58 netRa58 netL58 -3.0034432234306057e-13
Rbbr58 netL58 node_4 923.5928320471352
Cbr58 netL58 node_4 -4.1721648118982753e-19

* Branch 59
Rabr59 node_1 netRa59 373.4972256380368
Lbr59 netRa59 netL59 -6.580835750738872e-13
Rbbr59 netL59 node_4 -2764.8815430491263
Cbr59 netL59 node_4 -6.364795176250107e-19

* Branch 60
Rabr60 node_1 netRa60 70.45087793717506
Lbr60 netRa60 netL60 5.250283631578386e-13
Rbbr60 netL60 node_4 -1902.869258557501
Cbr60 netL60 node_4 3.9310460491248214e-18

* Branch 61
Rabr61 node_1 netRa61 1440.7136739490586
Lbr61 netRa61 netL61 2.7173121232902814e-12
Rbbr61 netL61 node_4 -3585.248855138147
Cbr61 netL61 node_4 5.265012536745596e-19

* Branch 62
Rabr62 node_1 netRa62 4078.40208604021
Lbr62 netRa62 netL62 1.7209946285846648e-11
Rbbr62 netL62 node_4 -58135.78323953897
Cbr62 netL62 node_4 7.2716242616548e-20

* Branch 63
Rabr63 node_1 netRa63 -32.072836082983876
Lbr63 netRa63 netL63 -2.9670746534975137e-13
Rbbr63 netL63 node_4 4269.412085211127
Cbr63 netL63 node_4 -2.17319125290927e-18

* Branch 64
Rabr64 node_1 netRa64 18.562767902588238
Lbr64 netRa64 netL64 2.1705159605682966e-12
Rbbr64 netL64 node_4 -203569.1374670802
Cbr64 netL64 node_4 5.95147953483225e-19

* Branch 65
Rabr65 node_1 netRa65 -1427.37801495402
Lbr65 netRa65 netL65 1.5036329573722688e-12
Rbbr65 netL65 node_4 2416.2421125420356
Cbr65 netL65 node_4 4.358439247827758e-19

* Branch 66
Rabr66 node_1 netRa66 -24523.146894329057
Lbr66 netRa66 netL66 2.2484544562965727e-11
Rbbr66 netL66 node_4 41131.891699456384
Cbr66 netL66 node_4 2.2286187555658893e-20

* Branch 67
Rabr67 node_1 netRa67 103222.35520496791
Lbr67 netRa67 netL67 -2.638138860148418e-11
Rbbr67 netL67 node_4 -108873.27702217131
Cbr67 netL67 node_4 -2.3473973102288122e-21

* Branch 68
Rabr68 node_1 netRa68 55.63559182151773
Lbr68 netRa68 netL68 -3.5669184237822286e-13
Rbbr68 netL68 node_4 -3676.7805926369488
Cbr68 netL68 node_4 -1.742709068293395e-18

* Branch 69
Rabr69 node_1 netRa69 5619.111195269547
Lbr69 netRa69 netL69 8.708802731390876e-12
Rbbr69 netL69 node_4 -17380.48400742838
Cbr69 netL69 node_4 8.918206286258471e-20

* Branch 70
Rabr70 node_1 netRa70 -852.6577828142163
Lbr70 netRa70 netL70 -8.493188420488771e-12
Rbbr70 netL70 node_4 34244.21583389086
Cbr70 netL70 node_4 -2.9089016426471343e-19

* Branch 71
Rabr71 node_1 netRa71 364.73730480256444
Lbr71 netRa71 netL71 -6.855043966287399e-13
Rbbr71 netL71 node_4 -2829.7396166605645
Cbr71 netL71 node_4 -6.641401501395658e-19

* Branch 72
Rabr72 node_1 netRa72 -2956.706179746978
Lbr72 netRa72 netL72 1.4177363849573107e-12
Rbbr72 netL72 node_4 3911.874746691965
Cbr72 netL72 node_4 1.2257145837846032e-19

* Branch 73
Rabr73 node_1 netRa73 -2709.691117179891
Lbr73 netRa73 netL73 -2.013487486323594e-12
Rbbr73 netL73 node_4 4876.96162717331
Cbr73 netL73 node_4 -1.523734881466803e-19

* Branch 74
Rabr74 node_1 netRa74 2383.4932328407017
Lbr74 netRa74 netL74 1.6970938228973755e-11
Rbbr74 netL74 node_4 -111877.32229349797
Cbr74 netL74 node_4 6.368952356149734e-20

* Branch 75
Rabr75 node_1 netRa75 640.7947315348663
Lbr75 netRa75 netL75 -3.2424877512529777e-12
Rbbr75 netL75 node_4 -27302.280118517974
Cbr75 netL75 node_4 -1.8521937690812447e-19

* Branch 76
Rabr76 node_1 netRa76 17.965750259215127
Lbr76 netRa76 netL76 1.2926291471613272e-12
Rbbr76 netL76 node_4 -64112.45934014199
Cbr76 netL76 node_4 1.1326066724338032e-18

* Branch 77
Rabr77 node_1 netRa77 -369.22006510788736
Lbr77 netRa77 netL77 -4.979662717093484e-13
Rbbr77 netL77 node_4 1371.6516594192603
Cbr77 netL77 node_4 -9.834489233761567e-19

* Branch 78
Rabr78 node_1 netRa78 -6673.234977602131
Lbr78 netRa78 netL78 5.305656792731508e-12
Rbbr78 netL78 node_4 13719.658173985872
Cbr78 netL78 node_4 5.794170263144011e-20

* Branch 79
Rabr79 node_1 netRa79 -326294.3830931333
Lbr79 netRa79 netL79 5.013417026969585e-11
Rbbr79 netL79 node_4 339524.42366981984
Cbr79 netL79 node_4 4.52520704328572e-22

* Branch 80
Rabr80 node_1 netRa80 -1790173.2697482847
Lbr80 netRa80 netL80 1.2873207678742739e-10
Rbbr80 netL80 node_4 1796215.8941098417
Cbr80 netL80 node_4 4.0033731574425795e-23

* Branch 81
Rabr81 node_1 netRa81 4815.710576142481
Lbr81 netRa81 netL81 1.593394205526572e-12
Rbbr81 netL81 node_4 -5386.617345606324
Cbr81 netL81 node_4 6.143008320165552e-20

* Branch 82
Rabr82 node_1 netRa82 -232978.42521793104
Lbr82 netRa82 netL82 -3.4760884977915704e-11
Rbbr82 netL82 node_4 242381.15002783158
Cbr82 netL82 node_4 -6.155908287182186e-22

* Branch 83
Rabr83 node_1 netRa83 1334.2808278890625
Lbr83 netRa83 netL83 2.5005099023789668e-12
Rbbr83 netL83 node_4 -5740.20939668496
Cbr83 netL83 node_4 3.2664115512554796e-19

* Branch 84
Rabr84 node_1 netRa84 -975.1073373259047
Lbr84 netRa84 netL84 -1.6325011477094276e-12
Rbbr84 netL84 node_4 5803.213348794753
Cbr84 netL84 node_4 -2.8862172938754764e-19

* Branch 85
Rabr85 node_1 netRa85 -1756.8976021061558
Lbr85 netRa85 netL85 -4.089881901988896e-12
Rbbr85 netL85 node_4 20441.498863221484
Cbr85 netL85 node_4 -1.1396235721699327e-19

* Branch 86
Rabr86 node_1 netRa86 -1590.2334659469777
Lbr86 netRa86 netL86 -1.8380030743221677e-12
Rbbr86 netL86 node_4 5548.517745557544
Cbr86 netL86 node_4 -2.0839509281732995e-19

* Branch 87
Rabr87 node_1 netRa87 95.83060500825106
Lbr87 netRa87 netL87 -1.314105202254343e-12
Rbbr87 netL87 node_4 -36178.49998894437
Cbr87 netL87 node_4 -3.770802190912131e-19

* Branch 88
Rabr88 node_1 netRa88 -5239.861026842191
Lbr88 netRa88 netL88 -2.7828400155822227e-12
Rbbr88 netL88 node_4 8365.104602791378
Cbr88 netL88 node_4 -6.350230674018197e-20

* Branch 89
Rabr89 node_1 netRa89 408.54238468405526
Lbr89 netRa89 netL89 2.6494016604176804e-12
Rbbr89 netL89 node_4 -18448.85310386966
Cbr89 netL89 node_4 3.5264434271027504e-19

* Branch 90
Rabr90 node_1 netRa90 -3341.041611291958
Lbr90 netRa90 netL90 -2.598157454111042e-12
Rbbr90 netL90 node_4 6095.886193073923
Cbr90 netL90 node_4 -1.2762123077430803e-19

* Branch 91
Rabr91 node_1 netRa91 4137.978925932567
Lbr91 netRa91 netL91 9.473307528524618e-12
Rbbr91 netL91 node_4 -25304.18706162924
Cbr91 netL91 node_4 9.05890077910592e-20

* Branch 92
Rabr92 node_1 netRa92 3507.5578659408807
Lbr92 netRa92 netL92 2.2181643353377624e-12
Rbbr92 netL92 node_4 -4925.74918097007
Cbr92 netL92 node_4 1.2843374518820048e-19

* Branch 93
Rabr93 node_1 netRa93 -321.88457902177663
Lbr93 netRa93 netL93 -9.59228428864707e-13
Rbbr93 netL93 node_4 6527.9246687381
Cbr93 netL93 node_4 -4.576968354243147e-19

* Branch 94
Rabr94 node_1 netRa94 -702.0733506015698
Lbr94 netRa94 netL94 -8.013867013713204e-13
Rbbr94 netL94 node_4 2731.228597235163
Cbr94 netL94 node_4 -4.183653540769606e-19

* Branch 95
Rabr95 node_1 netRa95 819.0942772566225
Lbr95 netRa95 netL95 -9.935925167625068e-13
Rbbr95 netL95 node_4 -3970.3396212849534
Cbr95 netL95 node_4 -3.046690242821169e-19

* Branch 96
Rabr96 node_1 netRa96 483.00494585064143
Lbr96 netRa96 netL96 1.4108780136194005e-13
Rbbr96 netL96 node_4 -596.4491207425353
Cbr96 netL96 node_4 4.909072685519903e-19

* Branch 97
Rabr97 node_1 netRa97 -67.0010354268781
Lbr97 netRa97 netL97 -2.0665664156821663e-13
Rbbr97 netL97 node_4 1750.7973042458514
Cbr97 netL97 node_4 -1.8755015018307156e-18

* Branch 98
Rabr98 node_1 netRa98 -53.408144363142924
Lbr98 netRa98 netL98 7.608853669882785e-14
Rbbr98 netL98 node_4 335.76660466938347
Cbr98 netL98 node_4 3.9130949593588766e-18

* Branch 99
Rabr99 node_1 netRa99 -5684.119792905749
Lbr99 netRa99 netL99 3.5863079086621333e-13
Rbbr99 netL99 node_4 5761.862501582405
Cbr99 netL99 node_4 1.0890496848464644e-20

.ends


* Y'22
.subckt yp22 node_2 0
* Branch 0
Rabr0 node_2 netRa0 -103541.61140550218
Lbr0 netRa0 netL0 -2.2500589839462288e-10
Rbbr0 netL0 0 1772231.900056806
Cbr0 netL0 0 -1.313621339499569e-21

* Branch 1
Rabr1 node_2 netRa1 -190304.8265284463
Lbr1 netRa1 netL1 -3.1863790930135565e-10
Rbbr1 netL1 0 1902762.347505642
Cbr1 netL1 0 -9.210451002306042e-22

* Branch 2
Rabr2 node_2 netRa2 -40004.72115537978
Lbr2 netRa2 netL2 -1.5177889724495803e-10
Rbbr2 netL2 0 2133689.1862066337
Cbr2 netL2 0 -1.9761581520084375e-21

* Branch 3
Rabr3 node_2 netRa3 -557900.3556684997
Lbr3 netRa3 netL3 -8.968955302974467e-10
Rbbr3 netL3 0 4103290.4671988506
Cbr3 netL3 0 -4.0657953665530313e-22

* Branch 4
Rabr4 node_2 netRa4 -437971.90970493923
Lbr4 netRa4 netL4 -6.884882560427238e-10
Rbbr4 netL4 0 3399403.719337138
Cbr4 netL4 0 -4.788291029897882e-22

* Branch 5
Rabr5 node_2 netRa5 -564570.3097605626
Lbr5 netRa5 netL5 -9.81046310848338e-10
Rbbr5 netL5 0 4560731.751271664
Cbr5 netL5 0 -3.9554733595346583e-22

* Branch 6
Rabr6 node_2 netRa6 -642277.3035732699
Lbr6 netRa6 netL6 -1.4049842637266513e-09
Rbbr6 netL6 0 6163211.712681353
Cbr6 netL6 0 -3.7184552341354247e-22

* Branch 7
Rabr7 node_2 netRa7 -499706.6042067385
Lbr7 netRa7 netL7 -7.74363968410906e-10
Rbbr7 netL7 0 3617142.7429275704
Cbr7 netL7 0 -4.421842836846314e-22

* Branch 8
Rabr8 node_2 netRa8 -645561.9555177588
Lbr8 netRa8 netL8 -1.324927400338113e-09
Rbbr8 netL8 0 5802059.960029343
Cbr8 netL8 0 -3.6863989403019787e-22

* Branch 9
Rabr9 node_2 netRa9 -641891.7618359991
Lbr9 netRa9 netL9 -1.5763762092192736e-09
Rbbr9 netL9 0 6789084.030242602
Cbr9 netL9 0 -3.7930694751807615e-22

* Branch 10
Rabr10 node_2 netRa10 -580751.2568245875
Lbr10 netRa10 netL10 -1.7930368432636782e-09
Rbbr10 netL10 0 7741749.93376096
Cbr10 netL10 0 -4.2125715790174813e-22

* Branch 11
Rabr11 node_2 netRa11 -622388.695048217
Lbr11 netRa11 netL11 -1.6587379875521932e-09
Rbbr11 netL11 0 7132610.377524151
Cbr11 netL11 0 -3.9157513047675483e-22

* Branch 12
Rabr12 node_2 netRa12 -433270.2253764261
Lbr12 netRa12 netL12 -1.9000833422155895e-09
Rbbr12 netL12 0 9779333.6892159
Cbr12 netL12 0 -4.814756394585634e-22

* Branch 13
Rabr13 node_2 netRa13 -541187.625580181
Lbr13 netRa13 netL13 -2.133755250147468e-09
Rbbr13 netL13 0 7814273.689789062
Cbr13 netL13 0 -5.360528943784755e-22

* Branch 14
Rabr14 node_2 netRa14 -577436.7888474601
Lbr14 netRa14 netL14 -6.25343989221591e-10
Rbbr14 netL14 0 2494578.2169828494
Cbr14 netL14 0 -4.409247070524292e-22

* Branch 15
Rabr15 node_2 netRa15 -406787.733613395
Lbr15 netRa15 netL15 -2.2830091155987967e-09
Rbbr15 netL15 0 8774510.680130411
Cbr15 netL15 0 -6.911401344834281e-22

* Branch 16
Rabr16 node_2 netRa16 -440052.372933752
Lbr16 netRa16 netL16 -2.2333868536203236e-09
Rbbr16 netL16 0 8562235.05735938
Cbr16 netL16 0 -6.330939703718819e-22

* Branch 17
Rabr17 node_2 netRa17 -616720.2296275228
Lbr17 netRa17 netL17 -1.153896996323038e-09
Rbbr17 netL17 0 5162848.593324174
Cbr17 netL17 0 -3.70759927756688e-22

* Branch 18
Rabr18 node_2 netRa18 -609085.2633804041
Lbr18 netRa18 netL18 -1.7256917677047691e-09
Rbbr18 netL18 0 7308211.580707376
Cbr18 netL18 0 -4.0054755096431824e-22

* Branch 19
Rabr19 node_2 netRa19 770727.9059850427
Lbr19 netRa19 netL19 -2.563208979502596e-10
Rbbr19 netL19 0 -1057162.798726317
Cbr19 netL19 0 -3.134098168764683e-22

* Branch 20
Rabr20 node_2 netRa20 -490237.34312950424
Lbr20 netRa20 netL20 -2.1804842265864315e-09
Rbbr20 netL20 0 8127381.25585693
Cbr20 netL20 0 -5.751636613890554e-22

* Branch 21
Rabr21 node_2 netRa21 -594001.6778723717
Lbr21 netRa21 netL21 -2.0695380685070744e-09
Rbbr21 netL21 0 7216273.369558624
Cbr21 netL21 0 -5.012209765366389e-22

* Branch 22
Rabr22 node_2 netRa22 -334668.47138512216
Lbr22 netRa22 netL22 -2.3810124278181797e-09
Rbbr22 netL22 0 9170733.654454963
Cbr22 netL22 0 -8.386524274688578e-22

* Branch 23
Rabr23 node_2 netRa23 -668912.430360645
Lbr23 netRa23 netL23 -1.2560500413551965e-09
Rbbr23 netL23 0 5307400.276303015
Cbr23 netL23 0 -3.60713581657389e-22

* Branch 24
Rabr24 node_2 netRa24 -31456.244323434676
Lbr24 netRa24 netL24 -5.072063356794042e-11
Rbbr24 netL24 0 321964.8852526384
Cbr24 netL24 0 -5.082220247477668e-21

* Branch 25
Rabr25 node_2 netRa25 -646996.5597837691
Lbr25 netRa25 netL25 -1.4909625721160706e-09
Rbbr25 netL25 0 6321771.744594099
Cbr25 netL25 0 -3.721818081086018e-22

* Branch 26
Rabr26 node_2 netRa26 -527983.1049644443
Lbr26 netRa26 netL26 -1.882921110184747e-09
Rbbr26 netL26 0 8329436.122289988
Cbr26 netL26 0 -4.406917318880424e-22

* Branch 27
Rabr27 node_2 netRa27 -377038.7645828149
Lbr27 netRa27 netL27 -2.3347199452995664e-09
Rbbr27 netL27 0 8627635.194057655
Cbr27 netL27 0 -7.525865951491111e-22

* Branch 28
Rabr28 node_2 netRa28 -841665.5657371221
Lbr28 netRa28 netL28 -1.9416671010823194e-09
Rbbr28 netL28 0 5184686.811790373
Cbr28 netL28 0 -4.524391808997395e-22

* Branch 29
Rabr29 node_2 netRa29 -251485.83800116507
Lbr29 netRa29 netL29 -3.0875102159538024e-10
Rbbr29 netL29 0 1366397.233746229
Cbr29 netL29 0 -9.064236229517817e-22

* Branch 30
Rabr30 node_2 netRa30 -669704.2844566343
Lbr30 netRa30 netL30 -1.1294113089020525e-09
Rbbr30 netL30 0 4670340.8762416765
Cbr30 netL30 0 -3.6251338570313086e-22

* Branch 31
Rabr31 node_2 netRa31 -6390833.874253104
Lbr31 netRa31 netL31 -1.017914314741712e-09
Rbbr31 netL31 0 6861771.584282749
Cbr31 netL31 0 -2.3219585480313093e-23

* Branch 32
Rabr32 node_2 netRa32 -561495.4904888683
Lbr32 netRa32 netL32 -1.8063737513419767e-10
Rbbr32 netL32 0 763936.9194532871
Cbr32 netL32 0 -4.2138543503740324e-22

* Branch 33
Rabr33 node_2 netRa33 192550.18237603075
Lbr33 netRa33 netL33 -6.293320702386951e-10
Rbbr33 netL33 0 -2191333.2828413458
Cbr33 netL33 0 -1.4850627193026479e-21

* Branch 34
Rabr34 node_2 netRa34 -289404.1397342406
Lbr34 netRa34 netL34 -1.6978483995782163e-10
Rbbr34 netL34 0 616964.8744023467
Cbr34 netL34 0 -9.513867992210049e-22

* Branch 35
Rabr35 node_2 netRa35 -284518.78575768403
Lbr35 netRa35 netL35 -9.287771479331275e-10
Rbbr35 netL35 0 7696644.689115099
Cbr35 netL35 0 -4.2502733914595915e-22

* Branch 36
Rabr36 node_2 netRa36 -401139.79793095874
Lbr36 netRa36 netL36 -5.316067336353925e-10
Rbbr36 netL36 0 2494806.687973439
Cbr36 netL36 0 -5.315549758864662e-22

* Branch 37
Rabr37 node_2 netRa37 -574045.9322263643
Lbr37 netRa37 netL37 -3.0218100226234455e-10
Rbbr37 netL37 0 1086751.3472048054
Cbr37 netL37 0 -4.844810232993564e-22

* Branch 38
Rabr38 node_2 netRa38 -711455.5522025183
Lbr38 netRa38 netL38 -4.0529867646182995e-10
Rbbr38 netL38 0 1440809.8807328246
Cbr38 netL38 0 -3.954510432562943e-22

* Branch 39
Rabr39 node_2 netRa39 -759260.3265078327
Lbr39 netRa39 netL39 -4.889686482378008e-10
Rbbr39 netL39 0 1733955.5130902643
Cbr39 netL39 0 -3.714708301853155e-22

* Branch 40
Rabr40 node_2 netRa40 -591840.1413771866
Lbr40 netRa40 netL40 -2.2934091530729884e-09
Rbbr40 netL40 0 8345449.794857978
Cbr40 netL40 0 -4.647924265043366e-22

* Branch 41
Rabr41 node_2 netRa41 -753689.0440190819
Lbr41 netRa41 netL41 -5.815391594140825e-10
Rbbr41 netL41 0 2114382.981116102
Cbr41 netL41 0 -3.649965504565167e-22

* Branch 42
Rabr42 node_2 netRa42 -782698.03876998
Lbr42 netRa42 netL42 -1.9731896253541166e-09
Rbbr42 netL42 0 9098148.103732623
Cbr42 netL42 0 -2.7723958059326807e-22

* Branch 43
Rabr43 node_2 netRa43 -158826.11530670736
Lbr43 netRa43 netL43 -3.1895364424696424e-09
Rbbr43 netL43 0 31683318.74379443
Cbr43 netL43 0 -6.36348587619258e-22

* Branch 44
Rabr44 node_2 netRa44 -1877916.7152345816
Lbr44 netRa44 netL44 -2.1205217718550645e-09
Rbbr44 netL44 0 4129201.0080916747
Cbr44 netL44 0 -2.735115895574937e-22

* Branch 45
Rabr45 node_2 netRa45 -1526670.466310708
Lbr45 netRa45 netL45 -1.468676398750953e-09
Rbbr45 netL45 0 4664063.574342513
Cbr45 netL45 0 -2.062894779031675e-22

* Branch 46
Rabr46 node_2 netRa46 -1379793.986601855
Lbr46 netRa46 netL46 -1.4762976514631787e-09
Rbbr46 netL46 0 4720333.81477277
Cbr46 netL46 0 -2.267009174620079e-22

* Branch 47
Rabr47 node_2 netRa47 -725464.848651993
Lbr47 netRa47 netL47 -3.122875507792049e-09
Rbbr47 netL47 0 9898252.908486148
Cbr47 netL47 0 -4.351296411683854e-22

* Branch 48
Rabr48 node_2 netRa48 -1991655.3550514034
Lbr48 netRa48 netL48 -9.519167216341458e-10
Rbbr48 netL48 0 3287275.8858449603
Cbr48 netL48 0 -1.454024399279176e-22

* Branch 49
Rabr49 node_2 netRa49 -807991.8988454824
Lbr49 netRa49 netL49 -4.147080007789875e-09
Rbbr49 netL49 0 15968640.316921167
Cbr49 netL49 0 -3.2158693085631695e-22

* Branch 50
Rabr50 node_2 netRa50 -730460.263904616
Lbr50 netRa50 netL50 -3.905441085515163e-09
Rbbr50 netL50 0 14364583.618073015
Cbr50 netL50 0 -3.7240965986748223e-22

* Branch 51
Rabr51 node_2 netRa51 -2053527.692112346
Lbr51 netRa51 netL51 -1.0172530677585595e-09
Rbbr51 netL51 0 3458158.1118031847
Cbr51 netL51 0 -1.432527525415974e-22

* Branch 52
Rabr52 node_2 netRa52 -472489.21852059977
Lbr52 netRa52 netL52 -5.356728093339058e-09
Rbbr52 netL52 0 28759216.055831637
Cbr52 netL52 0 -3.945926361096275e-22

* Branch 53
Rabr53 node_2 netRa53 -1922682.3827414361
Lbr53 netRa53 netL53 -1.2496617915327395e-09
Rbbr53 netL53 0 3996195.3563807546
Cbr53 netL53 0 -1.6265171734877278e-22

* Branch 54
Rabr54 node_2 netRa54 -1806656.9988144857
Lbr54 netRa54 netL54 -1.9199026446551414e-09
Rbbr54 netL54 0 5505736.640870669
Cbr54 netL54 0 -1.9302844988062617e-22

* Branch 55
Rabr55 node_2 netRa55 -2329125.9845079524
Lbr55 netRa55 netL55 -1.790850034275437e-09
Rbbr55 netL55 0 5765529.789696561
Cbr55 netL55 0 -1.3336764343372167e-22

* Branch 56
Rabr56 node_2 netRa56 -1665261.1206859883
Lbr56 netRa56 netL56 -2.411303759920875e-09
Rbbr56 netL56 0 4827088.983629224
Cbr56 netL56 0 -3.00003515291374e-22

* Branch 57
Rabr57 node_2 netRa57 -1811018.9201663963
Lbr57 netRa57 netL57 -1.5319892093053172e-09
Rbbr57 netL57 0 4619643.123614112
Cbr57 netL57 0 -1.8312538456308586e-22

* Branch 58
Rabr58 node_2 netRa58 -1897762.6671274751
Lbr58 netRa58 netL58 -1.93271050371569e-09
Rbbr58 netL58 0 5562090.615894087
Cbr58 netL58 0 -1.8311106120845542e-22

* Branch 59
Rabr59 node_2 netRa59 -1882926.7318248255
Lbr59 netRa59 netL59 -2.0381312508262586e-09
Rbbr59 netL59 0 5672243.373169945
Cbr59 netL59 0 -1.9084140252388988e-22

* Branch 60
Rabr60 node_2 netRa60 -1925693.3326475096
Lbr60 netRa60 netL60 -1.7726940002278124e-09
Rbbr60 netL60 0 5208220.73725335
Cbr60 netL60 0 -1.7675906063311599e-22

* Branch 61
Rabr61 node_2 netRa61 -872482.2492190985
Lbr61 netRa61 netL61 -3.6473735583974853e-09
Rbbr61 netL61 0 8736912.735553838
Cbr61 netL61 0 -4.78596522468216e-22

* Branch 62
Rabr62 node_2 netRa62 -1921616.2803559045
Lbr62 netRa62 netL62 -1.7927914066258588e-09
Rbbr62 netL62 0 5201457.9757612925
Cbr62 netL62 0 -1.7937355827762747e-22

* Branch 63
Rabr63 node_2 netRa63 -1630800.1839319058
Lbr63 netRa63 netL63 -2.664054841508344e-09
Rbbr63 netL63 0 7022806.093307534
Cbr63 netL63 0 -2.326293045614021e-22

* Branch 64
Rabr64 node_2 netRa64 -865927.691593436
Lbr64 netRa64 netL64 -4.325202345076269e-09
Rbbr64 netL64 0 10399069.126744458
Cbr64 netL64 0 -4.804264849778524e-22

* Branch 65
Rabr65 node_2 netRa65 -1598837.661107415
Lbr65 netRa65 netL65 -2.7211268199222707e-09
Rbbr65 netL65 0 7153168.663094827
Cbr65 netL65 0 -2.379443628042936e-22

* Branch 66
Rabr66 node_2 netRa66 -2125263.3798195263
Lbr66 netRa66 netL66 -1.442121370226659e-09
Rbbr66 netL66 0 4457801.215324756
Cbr66 netL66 0 -1.522213357786229e-22

* Branch 67
Rabr67 node_2 netRa67 -1475842.617219034
Lbr67 netRa67 netL67 -4.145934781593482e-09
Rbbr67 netL67 0 8742814.490665067
Cbr67 netL67 0 -3.2133686029648734e-22

* Branch 68
Rabr68 node_2 netRa68 -1304971.4769700451
Lbr68 netRa68 netL68 -4.126309434783416e-09
Rbbr68 netL68 0 8373643.6787273465
Cbr68 netL68 0 -3.776369903317869e-22

* Branch 69
Rabr69 node_2 netRa69 -3265168.140138044
Lbr69 netRa69 netL69 -3.797817330576787e-09
Rbbr69 netL69 0 10240576.617650358
Cbr69 netL69 0 -1.1358239015457195e-22

* Branch 70
Rabr70 node_2 netRa70 -6215914.007634336
Lbr70 netRa70 netL70 -1.3285144041782947e-08
Rbbr70 netL70 0 30017225.37177173
Cbr70 netL70 0 -7.120333766246703e-23

* Branch 71
Rabr71 node_2 netRa71 -2832214.4463050826
Lbr71 netRa71 netL71 -4.086277332700451e-09
Rbbr71 netL71 0 10373018.526844317
Cbr71 netL71 0 -1.3909050057431972e-22

* Branch 72
Rabr72 node_2 netRa72 -1354766.5102606458
Lbr72 netRa72 netL72 -4.004247449422511e-09
Rbbr72 netL72 0 8407182.223512927
Cbr72 netL72 0 -3.51566880517288e-22

* Branch 73
Rabr73 node_2 netRa73 -552972.5049512042
Lbr73 netRa73 netL73 -3.788230060120726e-09
Rbbr73 netL73 0 15307002.275373043
Cbr73 netL73 0 -4.475739361388526e-22

* Branch 74
Rabr74 node_2 netRa74 369851.95885948685
Lbr74 netRa74 netL74 -4.176939431504509e-09
Rbbr74 netL74 0 -20067951.98632948
Cbr74 netL74 0 -5.626610471233408e-22

* Branch 75
Rabr75 node_2 netRa75 -709008.0536046374
Lbr75 netRa75 netL75 -2.9772591704584247e-09
Rbbr75 netL75 0 18796952.884849254
Cbr75 netL75 0 -2.2342097422766125e-22

* Branch 76
Rabr76 node_2 netRa76 30762049.98735182
Lbr76 netRa76 netL76 -1.3956798015767608e-08
Rbbr76 netL76 0 -33261963.27099193
Cbr76 netL76 0 -1.3640102270930414e-23

* Branch 77
Rabr77 node_2 netRa77 -4338061.172462475
Lbr77 netRa77 netL77 -2.8476256042092006e-09
Rbbr77 netL77 0 6507701.637982404
Cbr77 netL77 0 -1.0087137728662351e-22

* Branch 78
Rabr78 node_2 netRa78 5235885.014381925
Lbr78 netRa78 netL78 -4.538645257235526e-09
Rbbr78 netL78 0 -9355308.085463088
Cbr78 netL78 0 -9.26544979876313e-23

* Branch 79
Rabr79 node_2 netRa79 1505374.1103155229
Lbr79 netRa79 netL79 -3.77014562232708e-09
Rbbr79 netL79 0 -11740772.83459333
Cbr79 netL79 0 -2.1329258512305047e-22

* Branch 80
Rabr80 node_2 netRa80 -3657920.7454734882
Lbr80 netRa80 netL80 2.9780956064941736e-09
Rbbr80 netL80 0 6959506.900102267
Cbr80 netL80 0 1.1697993064207742e-22

* Branch 81
Rabr81 node_2 netRa81 13458740.038858417
Lbr81 netRa81 netL81 5.259800481040313e-09
Rbbr81 netL81 0 -16344625.90673985
Cbr81 netL81 0 2.391101126061976e-23

* Branch 82
Rabr82 node_2 netRa82 1103588470.2354162
Lbr82 netRa82 netL82 6.037291868890788e-08
Rbbr82 netL82 0 -1106926515.6451387
Cbr82 netL82 0 4.9421666590238366e-26

* Branch 83
Rabr83 node_2 netRa83 69717105.84210823
Lbr83 netRa83 netL83 -1.7260250120355723e-08
Rbbr83 netL83 0 -72890096.1933184
Cbr83 netL83 0 -3.3965176960322834e-24

* Branch 84
Rabr84 node_2 netRa84 14524000.412938975
Lbr84 netRa84 netL84 7.74846138802218e-09
Rbbr84 netL84 0 -17722865.93711658
Cbr84 netL84 0 3.010284575875158e-23

* Branch 85
Rabr85 node_2 netRa85 504552808.942911
Lbr85 netRa85 netL85 4.451435374239294e-08
Rbbr85 netL85 0 -507717102.56285554
Cbr85 netL85 0 1.7376966557214374e-25

* Branch 86
Rabr86 node_2 netRa86 6287109.401517216
Lbr86 netRa86 netL86 -3.6576431926344314e-09
Rbbr86 netL86 0 -9743982.589044545
Cbr86 netL86 0 -5.970304893020492e-23

* Branch 87
Rabr87 node_2 netRa87 -680520.2537937723
Lbr87 netRa87 netL87 2.798232734702554e-09
Rbbr87 netL87 0 13585830.815766118
Cbr87 netL87 0 3.0256912360452453e-22

* Branch 88
Rabr88 node_2 netRa88 627073.5491554003
Lbr88 netRa88 netL88 1.7679785312528252e-09
Rbbr88 netL88 0 -9426635.57351613
Cbr88 netL88 0 2.991594108384828e-22

* Branch 89
Rabr89 node_2 netRa89 53817012.047772154
Lbr89 netRa89 netL89 1.2218624624692726e-08
Rbbr89 netL89 0 -57479181.45593845
Cbr89 netL89 0 3.950038344465184e-24

* Branch 90
Rabr90 node_2 netRa90 2975642.901064575
Lbr90 netRa90 netL90 3.0320203666386943e-09
Rbbr90 netL90 0 -7580354.191496801
Cbr90 netL90 0 1.344330288171755e-22

* Branch 91
Rabr91 node_2 netRa91 119070556.61200465
Lbr91 netRa91 netL91 -2.2005854789701928e-08
Rbbr91 netL91 0 -125310785.29824458
Cbr91 netL91 0 -1.4748137073512326e-24

* Branch 92
Rabr92 node_2 netRa92 2026163.9175827752
Lbr92 netRa92 netL92 2.0820782565602786e-09
Rbbr92 netL92 0 -6115169.289398238
Cbr92 netL92 0 1.6806214950570197e-22

* Branch 93
Rabr93 node_2 netRa93 419938.9262156866
Lbr93 netRa93 netL93 1.1453803201449783e-09
Rbbr93 netL93 0 -7527038.793742437
Cbr93 netL93 0 3.6248714200964737e-22

* Branch 94
Rabr94 node_2 netRa94 -50434.77202367509
Lbr94 netRa94 netL94 1.3384178076981853e-09
Rbbr94 netL94 0 73056437.11807463
Cbr94 netL94 0 3.619520493576473e-22

* Branch 95
Rabr95 node_2 netRa95 1104707.5538507162
Lbr95 netRa95 netL95 1.2604048944849522e-09
Rbbr95 netL95 0 -4453920.735505989
Cbr95 netL95 0 2.562063889896251e-22

* Branch 96
Rabr96 node_2 netRa96 -718061.0938388181
Lbr96 netRa96 netL96 7.662114904556774e-10
Rbbr96 netL96 0 2899983.205685799
Cbr96 netL96 0 3.678897082012463e-22

* Branch 97
Rabr97 node_2 netRa97 497379.5747852348
Lbr97 netRa97 netL97 8.82242007028575e-10
Rbbr97 netL97 0 -4584750.91624342
Cbr97 netL97 0 3.8705479178923674e-22

* Branch 98
Rabr98 node_2 netRa98 -1652894.1663094051
Lbr98 netRa98 netL98 7.633775751962333e-10
Rbbr98 netL98 0 2615093.4012180287
Cbr98 netL98 0 1.765758346282458e-22

* Branch 99
Rabr99 node_2 netRa99 -894978.0290387983
Lbr99 netRa99 netL99 2.530715189020535e-10
Rbbr99 netL99 0 1140156.277419157
Cbr99 netL99 0 2.4796520015635367e-22

.ends


* Y'23
.subckt yp23 node_2 node_3
* Branch 0
Rabr0 node_2 netRa0 -52.24748368418379
Lbr0 netRa0 netL0 7.68728346564235e-14
Rbbr0 netL0 node_3 400.2495872153511
Cbr0 netL0 node_3 3.263320094799024e-18

* Branch 1
Rabr1 node_2 netRa1 -38.721476515242266
Lbr1 netRa1 netL1 1.0906062575590872e-13
Rbbr1 netL1 node_3 901.6659384635273
Cbr1 netL1 node_3 2.535594510970064e-18

* Branch 2
Rabr2 node_2 netRa2 119947.79802025815
Lbr2 netRa2 netL2 2.747882659070191e-12
Rbbr2 netL2 node_3 -120165.85988941381
Cbr2 netL2 node_3 1.9096646532062095e-22

* Branch 3
Rabr3 node_2 netRa3 -62.988276778490246
Lbr3 netRa3 netL3 -3.6273046153255296e-14
Rbbr3 netL3 node_3 137.15820372936685
Cbr3 netL3 node_3 -4.354869677066534e-18

* Branch 4
Rabr4 node_2 netRa4 395.38842107890775
Lbr4 netRa4 netL4 -2.7272684975668903e-13
Rbbr4 netL4 node_3 -799.4432805405467
Cbr4 netL4 node_3 -8.373057615878151e-19

* Branch 5
Rabr5 node_2 netRa5 -819.3762851875132
Lbr5 netRa5 netL5 -5.111583419688877e-13
Rbbr5 netL5 node_3 1754.9627121596857
Cbr5 netL5 node_3 -3.6393963328212985e-19

* Branch 6
Rabr6 node_2 netRa6 67.56665305943356
Lbr6 netRa6 netL6 -1.2136658051951565e-13
Rbbr6 netL6 node_3 -641.0754495851864
Cbr6 netL6 node_3 -2.6286838688083044e-18

* Branch 7
Rabr7 node_2 netRa7 650.8120543625548
Lbr7 netRa7 netL7 -3.872258386540931e-13
Rbbr7 netL7 node_3 -1158.0910203674775
Cbr7 netL7 node_3 -5.029516362962946e-19

* Branch 8
Rabr8 node_2 netRa8 1343.0509192648003
Lbr8 netRa8 netL8 -7.436046901349257e-13
Rbbr8 netL8 node_3 -2497.3032394748707
Cbr8 netL8 node_3 -2.1745416582411543e-19

* Branch 9
Rabr9 node_2 netRa9 133.92936742421958
Lbr9 netRa9 netL9 -1.5370381722698404e-13
Rbbr9 netL9 node_3 -693.5813962929464
Cbr9 netL9 node_3 -1.5932903886391908e-18

* Branch 10
Rabr10 node_2 netRa10 291.55888991272667
Lbr10 netRa10 netL10 -1.8347933799176967e-13
Rbbr10 netL10 node_3 -612.8239792382503
Cbr10 netL10 node_3 -1.0058367570977864e-18

* Branch 11
Rabr11 node_2 netRa11 -849.6189447619222
Lbr11 netRa11 netL11 3.345989397788139e-13
Rbbr11 netL11 node_3 1223.085250319775
Cbr11 netL11 node_3 3.1794925877583494e-19

* Branch 12
Rabr12 node_2 netRa12 -487.3754573222147
Lbr12 netRa12 netL12 -3.4967785519502115e-13
Rbbr12 netL12 node_3 1299.2659907375157
Cbr12 netL12 node_3 -5.642971983997845e-19

* Branch 13
Rabr13 node_2 netRa13 63.75069318523818
Lbr13 netRa13 netL13 -2.1078920023960593e-13
Rbbr13 netL13 node_3 -751.7404863049304
Cbr13 netL13 node_3 -4.0906779433199635e-18

* Branch 14
Rabr14 node_2 netRa14 359.98574666116923
Lbr14 netRa14 netL14 -2.201137542156716e-13
Rbbr14 netL14 node_3 -687.8491803618367
Cbr14 netL14 node_3 -8.76878154181879e-19

* Branch 15
Rabr15 node_2 netRa15 64.66961594911463
Lbr15 netRa15 netL15 -1.8293969319058334e-13
Rbbr15 netL15 node_3 -939.7075760291722
Cbr15 netL15 node_3 -2.846340321885099e-18

* Branch 16
Rabr16 node_2 netRa16 743.7845006493274
Lbr16 netRa16 netL16 -3.0070198522612337e-13
Rbbr16 netL16 node_3 -1047.557137416389
Cbr16 netL16 node_3 -3.8288939356304123e-19

* Branch 17
Rabr17 node_2 netRa17 105.87870535839814
Lbr17 netRa17 netL17 -1.811839162040767e-13
Rbbr17 netL17 node_3 -685.167246491147
Cbr17 netL17 node_3 -2.4196040795610587e-18

* Branch 18
Rabr18 node_2 netRa18 -569.2797540148327
Lbr18 netRa18 netL18 -2.3086045315451516e-13
Rbbr18 netL18 node_3 828.0738985819739
Cbr18 netL18 node_3 -4.93415680324795e-19

* Branch 19
Rabr19 node_2 netRa19 51.59528475615802
Lbr19 netRa19 netL19 -1.8899705426697064e-13
Rbbr19 netL19 node_3 -1165.27302354709
Cbr19 netL19 node_3 -2.9490475564903177e-18

* Branch 20
Rabr20 node_2 netRa20 -1428.5250309968637
Lbr20 netRa20 netL20 -5.245626915055009e-13
Rbbr20 netL20 node_3 1870.7197086948229
Cbr20 netL20 node_3 -1.9752591016674962e-19

* Branch 21
Rabr21 node_2 netRa21 39.58186558524606
Lbr21 netRa21 netL21 -2.075915911073983e-13
Rbbr21 netL21 node_3 -1068.0190645779705
Cbr21 netL21 node_3 -4.512587316806811e-18

* Branch 22
Rabr22 node_2 netRa22 20.275962305566004
Lbr22 netRa22 netL22 -2.064069508890488e-13
Rbbr22 netL22 node_3 -2610.4954282825065
Cbr22 netL22 node_3 -3.3507025071199887e-18

* Branch 23
Rabr23 node_2 netRa23 2.4962554576018503
Lbr23 netRa23 netL23 -2.35307403440128e-13
Rbbr23 netL23 node_3 -7592.088176498783
Cbr23 netL23 node_3 -4.977614328211391e-18

* Branch 24
Rabr24 node_2 netRa24 -1712.5175635499638
Lbr24 netRa24 netL24 8.693576044175075e-13
Rbbr24 netL24 node_3 3005.6303178928993
Cbr24 netL24 node_3 1.676573128554764e-19

* Branch 25
Rabr25 node_2 netRa25 19.765814285777694
Lbr25 netRa25 netL25 -2.186216758343185e-13
Rbbr25 netL25 node_3 -2001.0017038712754
Cbr25 netL25 node_3 -4.779235851794294e-18

* Branch 26
Rabr26 node_2 netRa26 -51.51690097677509
Lbr26 netRa26 netL26 -3.1071845156138027e-13
Rbbr26 netL26 node_3 1344.4493305002543
Cbr26 netL26 node_3 -4.879764008980745e-18

* Branch 27
Rabr27 node_2 netRa27 -11774.59272070087
Lbr27 netRa27 netL27 1.3983718637808067e-12
Rbbr27 netL27 node_3 12241.37622402533
Cbr27 netL27 node_3 9.686671489382701e-21

* Branch 28
Rabr28 node_2 netRa28 13.940911221426271
Lbr28 netRa28 netL28 -2.159485641380206e-13
Rbbr28 netL28 node_3 -3973.1091016007526
Cbr28 netL28 node_3 -3.281427670162511e-18

* Branch 29
Rabr29 node_2 netRa29 -6.10942354513575
Lbr29 netRa29 netL29 -2.57544614832898e-13
Rbbr29 netL29 node_3 17178.47795809462
Cbr29 netL29 node_3 -4.985194766728719e-18

* Branch 30
Rabr30 node_2 netRa30 2006.2099166508083
Lbr30 netRa30 netL30 -1.1610853846328274e-12
Rbbr30 netL30 node_3 -4092.8517250104387
Cbr30 netL30 node_3 -1.4042944376432557e-19

* Branch 31
Rabr31 node_2 netRa31 -10841828.67390236
Lbr31 netRa31 netL31 9.881464419240313e-11
Rbbr31 netL31 node_3 10844552.35014799
Cbr31 netL31 node_3 8.40353797092447e-25

* Branch 32
Rabr32 node_2 netRa32 82.09870076807832
Lbr32 netRa32 netL32 -3.888498636649424e-13
Rbbr32 netL32 node_3 -1011.1923133882622
Cbr32 netL32 node_3 -4.464423047568888e-18

* Branch 33
Rabr33 node_2 netRa33 -3965.234739640224
Lbr33 netRa33 netL33 -2.1606094680153092e-12
Rbbr33 netL33 node_3 5297.374668119247
Cbr33 netL33 node_3 -1.0341783380292461e-19

* Branch 34
Rabr34 node_2 netRa34 43.46176767822072
Lbr34 netRa34 netL34 -2.0099950605654568e-13
Rbbr34 netL34 node_3 -1482.10753635232
Cbr34 netL34 node_3 -2.9886067562602686e-18

* Branch 35
Rabr35 node_2 netRa35 1858.7402372253848
Lbr35 netRa35 netL35 -9.814957962466577e-13
Rbbr35 netL35 node_3 -3614.1590079546872
Cbr35 netL35 node_3 -1.453869245336887e-19

* Branch 36
Rabr36 node_2 netRa36 169.43829331067252
Lbr36 netRa36 netL36 -1.8379261198290916e-13
Rbbr36 netL36 node_3 -580.1314073520663
Cbr36 netL36 node_3 -1.8523097623881003e-18

* Branch 37
Rabr37 node_2 netRa37 -113.80773867561517
Lbr37 netRa37 netL37 -3.5442635751654413e-13
Rbbr37 netL37 node_3 806.9464052439298
Cbr37 netL37 node_3 -3.9603428620341066e-18

* Branch 38
Rabr38 node_2 netRa38 -10.147735554302567
Lbr38 netRa38 netL38 -2.62874482228826e-13
Rbbr38 netL38 node_3 5870.986994473404
Cbr38 netL38 node_3 -5.473776791859745e-18

* Branch 39
Rabr39 node_2 netRa39 1562.6009641599373
Lbr39 netRa39 netL39 1.4890733318005527e-12
Rbbr39 netL39 node_3 -2379.744059334122
Cbr39 netL39 node_3 4.030844335496585e-19

* Branch 40
Rabr40 node_2 netRa40 -2318.1504555194692
Lbr40 netRa40 netL40 -3.0059667190815434e-12
Rbbr40 netL40 node_3 6918.625587377442
Cbr40 netL40 node_3 -1.8909935633238708e-19

* Branch 41
Rabr41 node_2 netRa41 -779.227426409283
Lbr41 netRa41 netL41 -8.969251871230823e-13
Rbbr41 netL41 node_3 4243.255839010631
Cbr41 netL41 node_3 -2.73384897083102e-19

* Branch 42
Rabr42 node_2 netRa42 -2469.5208294076465
Lbr42 netRa42 netL42 -2.7772618597901108e-12
Rbbr42 netL42 node_3 4192.093994503933
Cbr42 netL42 node_3 -2.700337806894982e-19

* Branch 43
Rabr43 node_2 netRa43 1051.1530419208816
Lbr43 netRa43 netL43 -1.0459860501618219e-12
Rbbr43 netL43 node_3 -2298.8973650491153
Cbr43 netL43 node_3 -4.3055648966173965e-19

* Branch 44
Rabr44 node_2 netRa44 73.29191628040465
Lbr44 netRa44 netL44 -1.9151492271295213e-13
Rbbr44 netL44 node_3 -320.4143761371799
Cbr44 netL44 node_3 -8.047835728874561e-18

* Branch 45
Rabr45 node_2 netRa45 888.6519094669763
Lbr45 netRa45 netL45 -6.366141365129184e-13
Rbbr45 netL45 node_3 -2127.300373131127
Cbr45 netL45 node_3 -3.3558555512827177e-19

* Branch 46
Rabr46 node_2 netRa46 158.52063242754005
Lbr46 netRa46 netL46 -5.891416159614604e-13
Rbbr46 netL46 node_3 -1437.3454721105102
Cbr46 netL46 node_3 -2.5527682982379886e-18

* Branch 47
Rabr47 node_2 netRa47 -66.60426264381611
Lbr47 netRa47 netL47 -3.200446189874763e-13
Rbbr47 netL47 node_3 2080.4989928471127
Cbr47 netL47 node_3 -2.346660947901045e-18

* Branch 48
Rabr48 node_2 netRa48 1196.486069100788
Lbr48 netRa48 netL48 1.3414284676611841e-12
Rbbr48 netL48 node_3 -3126.88461289509
Cbr48 netL48 node_3 3.592236396092835e-19

* Branch 49
Rabr49 node_2 netRa49 -4159.195880311193
Lbr49 netRa49 netL49 2.067690258522446e-12
Rbbr49 netL49 node_3 5397.3754890899
Cbr49 netL49 node_3 9.203096886140332e-20

* Branch 50
Rabr50 node_2 netRa50 3607.38566540998
Lbr50 netRa50 netL50 -2.5206744020563465e-12
Rbbr50 netL50 node_3 -8305.834831877735
Cbr50 netL50 node_3 -8.40467554261333e-20

* Branch 51
Rabr51 node_2 netRa51 593.8515022611434
Lbr51 netRa51 netL51 1.4199392283385784e-12
Rbbr51 netL51 node_3 -2265.394719750146
Cbr51 netL51 node_3 1.0589623252186664e-18

* Branch 52
Rabr52 node_2 netRa52 1961.9385101475818
Lbr52 netRa52 netL52 -1.700104795656478e-12
Rbbr52 netL52 node_3 -5807.4594934958495
Cbr52 netL52 node_3 -1.4904250505707504e-19

* Branch 53
Rabr53 node_2 netRa53 -6040.676079647535
Lbr53 netRa53 netL53 5.517363106738895e-12
Rbbr53 netL53 node_3 11493.784128593683
Cbr53 netL53 node_3 7.93851264353852e-20

* Branch 54
Rabr54 node_2 netRa54 714.0104498494087
Lbr54 netRa54 netL54 -1.0268063527413566e-12
Rbbr54 netL54 node_3 -4484.267325014882
Cbr54 netL54 node_3 -3.2024729801759953e-19

* Branch 55
Rabr55 node_2 netRa55 5128.658027481505
Lbr55 netRa55 netL55 7.029261652438307e-12
Rbbr55 netL55 node_3 -9389.905444592616
Cbr55 netL55 node_3 1.461576811380534e-19

* Branch 56
Rabr56 node_2 netRa56 1311.0039450500465
Lbr56 netRa56 netL56 3.8617148507183875e-12
Rbbr56 netL56 node_3 -19340.812622371057
Cbr56 netL56 node_3 1.5271080503626595e-19

* Branch 57
Rabr57 node_2 netRa57 2374.736050360193
Lbr57 netRa57 netL57 5.1347159117485636e-12
Rbbr57 netL57 node_3 -7554.908805958739
Cbr57 netL57 node_3 2.866446408833641e-19

* Branch 58
Rabr58 node_2 netRa58 263465.72542508197
Lbr58 netRa58 netL58 6.709423997259515e-11
Rbbr58 netL58 node_3 -270605.0424322171
Cbr58 netL58 node_3 9.412238600510975e-22

* Branch 59
Rabr59 node_2 netRa59 205283.10520329766
Lbr59 netRa59 netL59 7.264486329543173e-11
Rbbr59 netL59 node_3 -224380.10315213288
Cbr59 netL59 node_3 1.5774173509336727e-21

* Branch 60
Rabr60 node_2 netRa60 -69319.76039587625
Lbr60 netRa60 netL60 -3.774753006254364e-11
Rbbr60 netL60 node_3 83969.13101519008
Cbr60 netL60 node_3 -6.4867046931499555e-21

* Branch 61
Rabr61 node_2 netRa61 11332.76411321029
Lbr61 netRa61 netL61 1.2882200247153565e-11
Rbbr61 netL61 node_3 -22668.56514228241
Cbr61 netL61 node_3 5.016599137746216e-20

* Branch 62
Rabr62 node_2 netRa62 2486.5653879999877
Lbr62 netRa62 netL62 3.4159681199511884e-11
Rbbr62 netL62 node_3 -726475.947356964
Cbr62 netL62 node_3 1.899731871903125e-20

* Branch 63
Rabr63 node_2 netRa63 22755039.27127047
Lbr63 netRa63 netL63 1.5824013875305555e-09
Rbbr63 netL63 node_3 -22843690.47757394
Cbr63 netL63 node_3 3.0442592697917692e-24

* Branch 64
Rabr64 node_2 netRa64 -1907.6898710747105
Lbr64 netRa64 netL64 1.463257344916935e-11
Rbbr64 netL64 node_3 71823.72635570675
Cbr64 netL64 node_3 1.0658275670879965e-19

* Branch 65
Rabr65 node_2 netRa65 4179.37074713252
Lbr65 netRa65 netL65 -1.9101647827824913e-11
Rbbr65 netL65 node_3 -38601.71741067367
Cbr65 netL65 node_3 -1.1829406323615356e-19

* Branch 66
Rabr66 node_2 netRa66 35193.15735144438
Lbr66 netRa66 netL66 -2.7716641715244078e-11
Rbbr66 netL66 node_3 -53483.820106453975
Cbr66 netL66 node_3 -1.4723327589746003e-20

* Branch 67
Rabr67 node_2 netRa67 -2696.975075262678
Lbr67 netRa67 netL67 2.7584927893404538e-11
Rbbr67 netL67 node_3 584110.753720688
Cbr67 netL67 node_3 1.7493439806824774e-20

* Branch 68
Rabr68 node_2 netRa68 21691.97592867581
Lbr68 netRa68 netL68 1.3342420536454215e-11
Rbbr68 netL68 node_3 -30280.590928065158
Cbr68 netL68 node_3 2.0313267829536026e-20

* Branch 69
Rabr69 node_2 netRa69 230543.70486796353
Lbr69 netRa69 netL69 1.0807317474540796e-10
Rbbr69 netL69 node_3 -274678.56751620764
Cbr69 netL69 node_3 1.706655921583736e-21

* Branch 70
Rabr70 node_2 netRa70 -26525.217205412864
Lbr70 netRa70 netL70 -1.4120168666585001e-11
Rbbr70 netL70 node_3 38740.75507972134
Cbr70 netL70 node_3 -1.374093069345508e-20

* Branch 71
Rabr71 node_2 netRa71 -12259.85303760084
Lbr71 netRa71 netL71 -1.056994541949423e-11
Rbbr71 netL71 node_3 25449.31346752245
Cbr71 netL71 node_3 -3.387755741434676e-20

* Branch 72
Rabr72 node_2 netRa72 16913.549817167917
Lbr72 netRa72 netL72 -4.2046590237617566e-11
Rbbr72 netL72 node_3 -191485.679001114
Cbr72 netL72 node_3 -1.2980755794665568e-20

* Branch 73
Rabr73 node_2 netRa73 -20759.160992380996
Lbr73 netRa73 netL73 -6.356678697259135e-11
Rbbr73 netL73 node_3 310952.9610448743
Cbr73 netL73 node_3 -9.849296622207994e-21

* Branch 74
Rabr74 node_2 netRa74 -438953.62525541557
Lbr74 netRa74 netL74 6.12542358529177e-11
Rbbr74 netL74 node_3 455292.002124912
Cbr74 netL74 node_3 3.064946737468394e-22

* Branch 75
Rabr75 node_2 netRa75 30984.63917637481
Lbr75 netRa75 netL75 -4.310892055196723e-11
Rbbr75 netL75 node_3 -85263.37267071193
Cbr75 netL75 node_3 -1.6315387398963972e-20

* Branch 76
Rabr76 node_2 netRa76 78516054413.44095
Lbr76 netRa76 netL76 -1.0153442890335912e-07
Rbbr76 netL76 node_3 -78516140092.08604
Cbr76 netL76 node_3 -1.6470085880867288e-29

* Branch 77
Rabr77 node_2 netRa77 123.29197298163858
Lbr77 netRa77 netL77 1.1086906657422001e-11
Rbbr77 netL77 node_3 -687291.3507697097
Cbr77 netL77 node_3 1.3218435112930629e-19

* Branch 78
Rabr78 node_2 netRa78 138320.6339886877
Lbr78 netRa78 netL78 -3.7624010665502846e-11
Rbbr78 netL78 node_3 -147935.27324151195
Cbr78 netL78 node_3 -1.838606333461365e-21

* Branch 79
Rabr79 node_2 netRa79 19371.32060342955
Lbr79 netRa79 netL79 2.97965900359013e-11
Rbbr79 netL79 node_3 -100278.66653192633
Cbr79 netL79 node_3 1.5343823174429697e-20

* Branch 80
Rabr80 node_2 netRa80 -3471.7532609784375
Lbr80 netRa80 netL80 -3.977692669789725e-12
Rbbr80 netL80 node_3 14855.58245078635
Cbr80 netL80 node_3 -7.714370017067384e-20

* Branch 81
Rabr81 node_2 netRa81 -2921.2992157395906
Lbr81 netRa81 netL81 6.585508320420764e-12
Rbbr81 netL81 node_3 23757.527433305007
Cbr81 netL81 node_3 9.484083490015323e-20

* Branch 82
Rabr82 node_2 netRa82 21658.677057396162
Lbr82 netRa82 netL82 1.566069033742242e-11
Rbbr82 netL82 node_3 -41106.19738301166
Cbr82 netL82 node_3 1.7593197780658166e-20

* Branch 83
Rabr83 node_2 netRa83 -3983.41462249398
Lbr83 netRa83 netL83 1.2349092743098051e-11
Rbbr83 netL83 node_3 73311.91073870326
Cbr83 netL83 node_3 4.225326710532196e-20

* Branch 84
Rabr84 node_2 netRa84 503921036.4685008
Lbr84 netRa84 netL84 3.548396437069331e-09
Rbbr84 netL84 node_3 -503945387.3642005
Cbr84 netL84 node_3 1.39729194607891e-26

* Branch 85
Rabr85 node_2 netRa85 1124479.8356536264
Lbr85 netRa85 netL85 -9.472569282341419e-11
Rbbr85 netL85 node_3 -1132541.8327306246
Cbr85 netL85 node_3 -7.437894318316666e-23

* Branch 86
Rabr86 node_2 netRa86 6475.584940448752
Lbr86 netRa86 netL86 1.180193913088372e-11
Rbbr86 netL86 node_3 -33167.0135605046
Cbr86 netL86 node_3 5.498410952047815e-20

* Branch 87
Rabr87 node_2 netRa87 -40918.35266537568
Lbr87 netRa87 netL87 1.037781544653578e-10
Rbbr87 netL87 node_3 530404.9599259344
Cbr87 netL87 node_3 4.7773751388956515e-21

* Branch 88
Rabr88 node_2 netRa88 -513.0658972918366
Lbr88 netRa88 netL88 -2.1495333286516934e-12
Rbbr88 netL88 node_3 21567.9429979336
Cbr88 netL88 node_3 -1.9456918559931058e-19

* Branch 89
Rabr89 node_2 netRa89 2108.8558906783423
Lbr89 netRa89 netL89 5.823183495307453e-12
Rbbr89 netL89 node_3 -24039.20207899808
Cbr89 netL89 node_3 1.1500109018406233e-19

* Branch 90
Rabr90 node_2 netRa90 2485.8036981598957
Lbr90 netRa90 netL90 1.6575296489568398e-11
Rbbr90 netL90 node_3 -148940.3930378966
Cbr90 netL90 node_3 4.48966405278588e-20

* Branch 91
Rabr91 node_2 netRa91 422280.3536367095
Lbr91 netRa91 netL91 2.578520699786589e-10
Rbbr91 netL91 node_3 -739030.09969854
Cbr91 netL91 node_3 8.264641671731532e-22

* Branch 92
Rabr92 node_2 netRa92 -21570.27282744295
Lbr92 netRa92 netL92 -1.542014254279104e-11
Rbbr92 netL92 node_3 45457.32432142397
Cbr92 netL92 node_3 -1.5732411779774512e-20

* Branch 93
Rabr93 node_2 netRa93 -37661.67784249955
Lbr93 netRa93 netL93 1.9297446766365935e-11
Rbbr93 netL93 node_3 57040.13225256047
Cbr93 netL93 node_3 8.98048582233341e-21

* Branch 94
Rabr94 node_2 netRa94 -229418.30405611818
Lbr94 netRa94 netL94 2.708791611754621e-11
Rbbr94 netL94 node_3 236177.59616818302
Cbr94 netL94 node_3 4.998918235045023e-22

* Branch 95
Rabr95 node_2 netRa95 -163.89542120891164
Lbr95 netRa95 netL95 9.158221698020135e-12
Rbbr95 netL95 node_3 1204240.4651826096
Cbr95 netL95 node_3 4.474844895959364e-20

* Branch 96
Rabr96 node_2 netRa96 -1875175.618487941
Lbr96 netRa96 netL96 1.4211402068459795e-10
Rbbr96 netL96 node_3 1900872.999875675
Cbr96 netL96 node_3 3.9867218143681966e-23

* Branch 97
Rabr97 node_2 netRa97 -20305.64129879382
Lbr97 netRa97 netL97 1.1093941689112143e-11
Rbbr97 netL97 node_3 33740.911853956546
Cbr97 netL97 node_3 1.6181378203105182e-20

* Branch 98
Rabr98 node_2 netRa98 -4161.851052933084
Lbr98 netRa98 netL98 4.811877571610268e-13
Rbbr98 netL98 node_3 4321.350052310023
Cbr98 netL98 node_3 2.6656729365073078e-20

* Branch 99
Rabr99 node_2 netRa99 -32.76810897611458
Lbr99 netRa99 netL99 5.236665068807964e-14
Rbbr99 netL99 node_3 288.0803257668642
Cbr99 netL99 node_3 4.8678418260232924e-18

.ends


* Y'24
.subckt yp24 node_2 node_4
* Branch 0
Rabr0 node_2 netRa0 11.496715003528813
Lbr0 netRa0 netL0 -2.1921305987062518e-14
Rbbr0 netL0 node_4 -112.99536336717546
Cbr0 netL0 node_4 -1.4641562994846602e-17

* Branch 1
Rabr1 node_2 netRa1 3.4535531046191146
Lbr1 netRa1 netL1 -2.646386305902219e-14
Rbbr1 netL1 node_4 -373.53176388274545
Cbr1 netL1 node_4 -1.336073464131234e-17

* Branch 2
Rabr2 node_2 netRa2 10.01804798818773
Lbr2 netRa2 netL2 -4.422855459798514e-14
Rbbr2 netL2 node_4 -536.9765748540738
Cbr2 netL2 node_4 -6.459764900328478e-18

* Branch 3
Rabr3 node_2 netRa3 -770.076523243319
Lbr3 netRa3 netL3 -1.3387100049702896e-13
Rbbr3 netL3 node_4 850.9050688195501
Cbr3 netL3 node_4 -2.064738557155289e-19

* Branch 4
Rabr4 node_2 netRa4 -2.1243245496851553
Lbr4 netRa4 netL4 1.8506017798356205e-14
Rbbr4 netL4 node_4 370.2775035361198
Cbr4 netL4 node_4 1.5647409984926144e-17

* Branch 5
Rabr5 node_2 netRa5 -37.93884674358672
Lbr5 netRa5 netL5 -5.279341052769202e-14
Rbbr5 netL5 node_4 261.68384502662013
Cbr5 netL5 node_4 -5.780272580558638e-18

* Branch 6
Rabr6 node_2 netRa6 -292.52310104850926
Lbr6 netRa6 netL6 -7.327696275338937e-14
Rbbr6 netL6 node_4 344.8727391965627
Cbr6 netL6 node_4 -7.358361730213205e-19

* Branch 7
Rabr7 node_2 netRa7 1080.6428930277953
Lbr7 netRa7 netL7 -2.4875015238378615e-13
Rbbr7 netL7 node_4 -1206.8755767141474
Cbr7 netL7 node_4 -1.888529436059995e-19

* Branch 8
Rabr8 node_2 netRa8 -63.465288882242504
Lbr8 netRa8 netL8 -4.946859209156838e-14
Rbbr8 netL8 node_4 196.67648130460537
Cbr8 netL8 node_4 -4.098259071508581e-18

* Branch 9
Rabr9 node_2 netRa9 -28.36139416137223
Lbr9 netRa9 netL9 2.5790028960850185e-14
Rbbr9 netL9 node_4 92.10579226768535
Cbr9 netL9 node_4 9.55659893027689e-18

* Branch 10
Rabr10 node_2 netRa10 385.84594087933687
Lbr10 netRa10 netL10 -1.0022342706158479e-13
Rbbr10 netL10 node_4 -444.423555644368
Cbr10 netL10 node_4 -5.79119865389631e-19

* Branch 11
Rabr11 node_2 netRa11 41.53856182168547
Lbr11 netRa11 netL11 2.9914747618259914e-14
Rbbr11 netL11 node_4 -102.68038557092767
Cbr11 netL11 node_4 7.174372110666947e-18

* Branch 12
Rabr12 node_2 netRa12 4039.04564009329
Lbr12 netRa12 netL12 5.158264832439096e-13
Rbbr12 netL12 node_4 -4194.75162588437
Cbr12 netL12 node_4 3.0565868899093733e-20

* Branch 13
Rabr13 node_2 netRa13 4.781666201073042
Lbr13 netRa13 netL13 -3.3211124678910435e-14
Rbbr13 netL13 node_4 -477.46548021623744
Cbr13 netL13 node_4 -1.2011331283015665e-17

* Branch 14
Rabr14 node_2 netRa14 -142097988.39708787
Lbr14 netRa14 netL14 -1.160228395322078e-10
Rbbr14 netL14 node_4 142098278.78898177
Cbr14 netL14 node_4 -5.7461404705077245e-27

* Branch 15
Rabr15 node_2 netRa15 6.60204266637173
Lbr15 netRa15 netL15 -2.116597868701992e-14
Rbbr15 netL15 node_4 -165.02597023748663
Cbr15 netL15 node_4 -1.7920896752356836e-17

* Branch 16
Rabr16 node_2 netRa16 -47419.54438176855
Lbr16 netRa16 netL16 -2.419401503002016e-12
Rbbr16 netL16 node_4 47789.83023789784
Cbr16 netL16 node_4 -1.0687471148043678e-21

* Branch 17
Rabr17 node_2 netRa17 -1027.8418027433377
Lbr17 netRa17 netL17 3.3188509736141286e-13
Rbbr17 netL17 node_4 1338.7226262969316
Cbr17 netL17 node_4 2.396280352434038e-19

* Branch 18
Rabr18 node_2 netRa18 67.85238628647643
Lbr18 netRa18 netL18 4.6258500666478433e-14
Rbbr18 netL18 node_4 -126.41681815560936
Cbr18 netL18 node_4 5.464784443610319e-18

* Branch 19
Rabr19 node_2 netRa19 28.48053102000418
Lbr19 netRa19 netL19 3.5008265961851675e-14
Rbbr19 netL19 node_4 -75.88038124711622
Cbr19 netL19 node_4 1.6574002169497588e-17

* Branch 20
Rabr20 node_2 netRa20 78.4466823846394
Lbr20 netRa20 netL20 4.9243569913978664e-14
Rbbr20 netL20 node_4 -132.29716436902282
Cbr20 netL20 node_4 4.7986320058589915e-18

* Branch 21
Rabr21 node_2 netRa21 -1407.3258044567028
Lbr21 netRa21 netL21 4.3785076214747776e-13
Rbbr21 netL21 node_4 1867.6743448134255
Cbr21 netL21 node_4 1.6568528529498198e-19

* Branch 22
Rabr22 node_2 netRa22 58.62980281602229
Lbr22 netRa22 netL22 4.743959640119161e-14
Rbbr22 netL22 node_4 -134.21707810913026
Cbr22 netL22 node_4 6.1092153645350535e-18

* Branch 23
Rabr23 node_2 netRa23 69.64902527207086
Lbr23 netRa23 netL23 5.924080993606703e-14
Rbbr23 netL23 node_4 -113.32667048117027
Cbr23 netL23 node_4 7.61076403704016e-18

* Branch 24
Rabr24 node_2 netRa24 89.5213650555781
Lbr24 netRa24 netL24 5.515583063241099e-14
Rbbr24 netL24 node_4 -139.55934573700458
Cbr24 netL24 node_4 4.459050820388002e-18

* Branch 25
Rabr25 node_2 netRa25 53.72329628840581
Lbr25 netRa25 netL25 6.177721826518849e-14
Rbbr25 netL25 node_4 -205.61471175786025
Cbr25 netL25 node_4 5.691722261929606e-18

* Branch 26
Rabr26 node_2 netRa26 -3468.1037980630053
Lbr26 netRa26 netL26 9.033890828132513e-13
Rbbr26 netL26 node_4 4100.160063433116
Cbr26 netL26 node_4 6.329764070046122e-20

* Branch 27
Rabr27 node_2 netRa27 59.86139886352994
Lbr27 netRa27 netL27 5.221988489557056e-14
Rbbr27 netL27 node_4 -103.39605384085527
Cbr27 netL27 node_4 8.53613538392932e-18

* Branch 28
Rabr28 node_2 netRa28 170202.31468860537
Lbr28 netRa28 netL28 3.705712267828174e-12
Rbbr28 netL28 node_4 -170293.61602431067
Cbr28 netL28 node_4 1.2788905825237096e-22

* Branch 29
Rabr29 node_2 netRa29 -6961.619814741594
Lbr29 netRa29 netL29 1.659293215757751e-12
Rbbr29 netL29 node_4 8195.480434772531
Cbr29 netL29 node_4 2.899489847420613e-20

* Branch 30
Rabr30 node_2 netRa30 79.15103607000903
Lbr30 netRa30 netL30 6.74183135470948e-14
Rbbr30 netL30 node_4 -124.47853594207814
Cbr30 netL30 node_4 6.91595800683063e-18

* Branch 31
Rabr31 node_2 netRa31 44.41740399716209
Lbr31 netRa31 netL31 4.293599516387522e-14
Rbbr31 netL31 node_4 -87.73817311610475
Cbr31 netL31 node_4 1.1150940527501609e-17

* Branch 32
Rabr32 node_2 netRa32 24449.005369819035
Lbr32 netRa32 netL32 -2.480424518276254e-12
Rbbr32 netL32 node_4 -25267.25030012004
Cbr32 netL32 node_4 -4.010611140706794e-21

* Branch 33
Rabr33 node_2 netRa33 134.92302601579286
Lbr33 netRa33 netL33 1.0018323998678999e-13
Rbbr33 netL33 node_4 -182.51662452050985
Cbr33 netL33 node_4 4.099319040178797e-18

* Branch 34
Rabr34 node_2 netRa34 83.41462794538016
Lbr34 netRa34 netL34 5.3406033448648185e-14
Rbbr34 netL34 node_4 -139.61975616433742
Cbr34 netL34 node_4 4.6155282188478885e-18

* Branch 35
Rabr35 node_2 netRa35 -3163.598011308006
Lbr35 netRa35 netL35 8.140925515557284e-13
Rbbr35 netL35 node_4 3709.0967571097995
Cbr35 netL35 node_4 6.921612131878784e-20

* Branch 36
Rabr36 node_2 netRa36 84.28403135119527
Lbr36 netRa36 netL36 5.441638277973524e-14
Rbbr36 netL36 node_4 -133.56281443668854
Cbr36 netL36 node_4 4.859529725688289e-18

* Branch 37
Rabr37 node_2 netRa37 32.08087521144903
Lbr37 netRa37 netL37 7.22403267473396e-14
Rbbr37 netL37 node_4 -119.69247125918672
Cbr37 netL37 node_4 1.9157538868840274e-17

* Branch 38
Rabr38 node_2 netRa38 84.39071820626829
Lbr38 netRa38 netL38 7.31829273611108e-14
Rbbr38 netL38 node_4 -129.03081399977077
Cbr38 netL38 node_4 6.766081912628104e-18

* Branch 39
Rabr39 node_2 netRa39 -185.2506157702137
Lbr39 netRa39 netL39 2.101072565969e-13
Rbbr39 netL39 node_4 320.54302639314017
Cbr39 netL39 node_4 3.5095917473150156e-18

* Branch 40
Rabr40 node_2 netRa40 303.45383232483744
Lbr40 netRa40 netL40 3.5770116385645023e-13
Rbbr40 netL40 node_4 -536.5645931736117
Cbr40 netL40 node_4 2.21413300415762e-18

* Branch 41
Rabr41 node_2 netRa41 2729.9229742010157
Lbr41 netRa41 netL41 7.486750962511462e-13
Rbbr41 netL41 node_4 -2971.4411469140014
Cbr41 netL41 node_4 9.245613037381733e-20

* Branch 42
Rabr42 node_2 netRa42 408.18749607249134
Lbr42 netRa42 netL42 1.7529105521113886e-13
Rbbr42 netL42 node_4 -454.1940949624562
Cbr42 netL42 node_4 9.475298152758757e-19

* Branch 43
Rabr43 node_2 netRa43 8.788795562970936
Lbr43 netRa43 netL43 2.960863932409669e-14
Rbbr43 netL43 node_4 -59.65178912325344
Cbr43 netL43 node_4 5.742934659318103e-17

* Branch 44
Rabr44 node_2 netRa44 116.31573221025882
Lbr44 netRa44 netL44 6.583752435448217e-14
Rbbr44 netL44 node_4 -165.02624382471754
Cbr44 netL44 node_4 3.4394935382772997e-18

* Branch 45
Rabr45 node_2 netRa45 494.37787240676096
Lbr45 netRa45 netL45 1.6589183157833533e-13
Rbbr45 netL45 node_4 -562.1375745888698
Cbr45 netL45 node_4 5.977578901298387e-19

* Branch 46
Rabr46 node_2 netRa46 47.393565353979504
Lbr46 netRa46 netL46 1.269463270140327e-13
Rbbr46 netL46 node_4 -251.05258049811982
Cbr46 netL46 node_4 1.0769041055657527e-17

* Branch 47
Rabr47 node_2 netRa47 9264.788309049916
Lbr47 netRa47 netL47 1.937360895875792e-12
Rbbr47 netL47 node_4 -10603.586025820248
Cbr47 netL47 node_4 1.9732566926204688e-20

* Branch 48
Rabr48 node_2 netRa48 -166976.91095155018
Lbr48 netRa48 netL48 4.6719373208033214e-12
Rbbr48 netL48 node_4 167311.29012385887
Cbr48 netL48 node_4 1.6721845142587151e-22

* Branch 49
Rabr49 node_2 netRa49 650.4987572153055
Lbr49 netRa49 netL49 2.6043363666132944e-13
Rbbr49 netL49 node_4 -895.916320039198
Cbr49 netL49 node_4 4.472116756676482e-19

* Branch 50
Rabr50 node_2 netRa50 -6394.046975746934
Lbr50 netRa50 netL50 -1.1319531110557865e-12
Rbbr50 netL50 node_4 6635.52463150507
Cbr50 netL50 node_4 -2.6687182222801387e-20

* Branch 51
Rabr51 node_2 netRa51 -3494.988501006946
Lbr51 netRa51 netL51 -1.1269620602043434e-12
Rbbr51 netL51 node_4 3888.475208523313
Cbr51 netL51 node_4 -8.294139662555724e-20

* Branch 52
Rabr52 node_2 netRa52 -1747.237152742379
Lbr52 netRa52 netL52 -7.536416256608963e-13
Rbbr52 netL52 node_4 2164.0683509938685
Cbr52 netL52 node_4 -1.993537709511059e-19

* Branch 53
Rabr53 node_2 netRa53 22441.01760034892
Lbr53 netRa53 netL53 -5.971621612763221e-12
Rbbr53 netL53 node_4 -23573.629391524657
Cbr53 netL53 node_4 -1.1287390516885517e-20

* Branch 54
Rabr54 node_2 netRa54 -497.55457975319626
Lbr54 netRa54 netL54 -7.017269676633636e-13
Rbbr54 netL54 node_4 983.2876737531168
Cbr54 netL54 node_4 -1.4348399701933388e-18

* Branch 55
Rabr55 node_2 netRa55 -5237.0252822653365
Lbr55 netRa55 netL55 -3.26513643779154e-12
Rbbr55 netL55 node_4 6136.2045188969105
Cbr55 netL55 node_4 -1.0161963950682126e-19

* Branch 56
Rabr56 node_2 netRa56 -52548.76198402009
Lbr56 netRa56 netL56 -1.6271892334121465e-11
Rbbr56 netL56 node_4 56292.198297910356
Cbr56 netL56 node_4 -5.501112892416828e-21

* Branch 57
Rabr57 node_2 netRa57 -1130.2010397152083
Lbr57 netRa57 netL57 -2.430840843358427e-12
Rbbr57 netL57 node_4 5177.745150053311
Cbr57 netL57 node_4 -4.154618452207846e-19

* Branch 58
Rabr58 node_2 netRa58 -577.4551035766997
Lbr58 netRa58 netL58 -2.2193866243417674e-12
Rbbr58 netL58 node_4 5904.564696113143
Cbr58 netL58 node_4 -6.510737405865966e-19

* Branch 59
Rabr59 node_2 netRa59 -8530.027080983595
Lbr59 netRa59 netL59 -9.541858494764928e-12
Rbbr59 netL59 node_4 12989.611183912959
Cbr59 netL59 node_4 -8.611720821054987e-20

* Branch 60
Rabr60 node_2 netRa60 -757.487530861882
Lbr60 netRa60 netL60 -1.2380176435977116e-12
Rbbr60 netL60 node_4 1700.1180194719975
Cbr60 netL60 node_4 -9.613447986634805e-19

* Branch 61
Rabr61 node_2 netRa61 -42242.49949293149
Lbr61 netRa61 netL61 -8.774483870538777e-11
Rbbr61 netL61 node_4 189109.9542541283
Cbr61 netL61 node_4 -1.0984547986695888e-20

* Branch 62
Rabr62 node_2 netRa62 4916.594966805757
Lbr62 netRa62 netL62 3.697498801579704e-12
Rbbr62 netL62 node_4 -10654.901723280824
Cbr62 netL62 node_4 7.058490938253922e-20

* Branch 63
Rabr63 node_2 netRa63 -265.7085306246773
Lbr63 netRa63 netL63 4.639055376429859e-12
Rbbr63 netL63 node_4 68067.39697881571
Cbr63 netL63 node_4 2.5618506920707343e-19

* Branch 64
Rabr64 node_2 netRa64 461.4196627969543
Lbr64 netRa64 netL64 3.934607376375578e-12
Rbbr64 netL64 node_4 -13724.53420582829
Cbr64 netL64 node_4 6.222880326603149e-19

* Branch 65
Rabr65 node_2 netRa65 -104819.34107203485
Lbr65 netRa65 netL65 -2.4674559224096555e-11
Rbbr65 netL65 node_4 109880.47967317984
Cbr65 netL65 node_4 -2.1424338048695105e-21

* Branch 66
Rabr66 node_2 netRa66 -442.5748982604928
Lbr66 netRa66 netL66 3.049561883978585e-13
Rbbr66 netL66 node_4 967.8895266744385
Cbr66 netL66 node_4 7.118117749720418e-19

* Branch 67
Rabr67 node_2 netRa67 -561.722468913874
Lbr67 netRa67 netL67 -1.6603508231922682e-11
Rbbr67 netL67 node_4 323091.77256718854
Cbr67 netL67 node_4 -9.21061899585374e-20

* Branch 68
Rabr68 node_2 netRa68 -3617.9118949307413
Lbr68 netRa68 netL68 -2.345084619550137e-12
Rbbr68 netL68 node_4 4655.581096876659
Cbr68 netL68 node_4 -1.3924897396530757e-19

* Branch 69
Rabr69 node_2 netRa69 -2584.063516863297
Lbr69 netRa69 netL69 -2.632735568518024e-12
Rbbr69 netL69 node_4 6240.089666539344
Cbr69 netL69 node_4 -1.633152457225735e-19

* Branch 70
Rabr70 node_2 netRa70 -228.90711062065776
Lbr70 netRa70 netL70 -6.584067769371231e-13
Rbbr70 netL70 node_4 3309.582776012278
Cbr70 netL70 node_4 -8.697495208607079e-19

* Branch 71
Rabr71 node_2 netRa71 -4749.056012260354
Lbr71 netRa71 netL71 -5.735078146640973e-12
Rbbr71 netL71 node_4 16323.005601407778
Cbr71 netL71 node_4 -7.40087138763551e-20

* Branch 72
Rabr72 node_2 netRa72 -53615.75193601224
Lbr72 netRa72 netL72 1.672569640383376e-11
Rbbr72 netL72 node_4 58339.38648965553
Cbr72 netL72 node_4 5.346740999316579e-21

* Branch 73
Rabr73 node_2 netRa73 -7908.391936473894
Lbr73 netRa73 netL73 -6.415922953408861e-12
Rbbr73 netL73 node_4 16141.229452867361
Cbr73 netL73 node_4 -5.027393485140223e-20

* Branch 74
Rabr74 node_2 netRa74 -905569.8233885174
Lbr74 netRa74 netL74 3.5313903696595706e-11
Rbbr74 netL74 node_4 906863.9417421309
Cbr74 netL74 node_4 4.3000747484454424e-23

* Branch 75
Rabr75 node_2 netRa75 280.44954892938495
Lbr75 netRa75 netL75 -8.242708061435628e-13
Rbbr75 netL75 node_4 -3784.1422866890302
Cbr75 netL75 node_4 -7.758693365855211e-19

* Branch 76
Rabr76 node_2 netRa76 11280.71456572749
Lbr76 netRa76 netL76 -3.5653967058120346e-12
Rbbr76 netL76 node_4 -13435.391338320213
Cbr76 netL76 node_4 -2.3521684028621212e-20

* Branch 77
Rabr77 node_2 netRa77 -4107.380730248429
Lbr77 netRa77 netL77 -2.5300882728480666e-12
Rbbr77 netL77 node_4 6784.6993928044485
Cbr77 netL77 node_4 -9.081252738041139e-20

* Branch 78
Rabr78 node_2 netRa78 -10794.431890496067
Lbr78 netRa78 netL78 -4.993841578584996e-12
Rbbr78 netL78 node_4 14983.353424888901
Cbr78 netL78 node_4 -3.0882088997122e-20

* Branch 79
Rabr79 node_2 netRa79 10954.661778855456
Lbr79 netRa79 netL79 3.35090591716808e-12
Rbbr79 netL79 node_4 -12529.717435207936
Cbr79 netL79 node_4 2.4416143373059372e-20

* Branch 80
Rabr80 node_2 netRa80 -24732.158715131376
Lbr80 netRa80 netL80 -4.848914321845695e-12
Rbbr80 netL80 node_4 25727.159219580688
Cbr80 netL80 node_4 -7.621265379663164e-21

* Branch 81
Rabr81 node_2 netRa81 156021.59700061468
Lbr81 netRa81 netL81 1.4569370980625246e-11
Rbbr81 netL81 node_4 -157710.14250487398
Cbr81 netL81 node_4 5.921298028764379e-22

* Branch 82
Rabr82 node_2 netRa82 -1067698.76575239
Lbr82 netRa82 netL82 -6.979454130839845e-11
Rbbr82 netL82 node_4 1072146.156974972
Cbr82 netL82 node_4 -6.097237934297378e-23

* Branch 83
Rabr83 node_2 netRa83 724.0002621092933
Lbr83 netRa83 netL83 -5.048876761597274e-13
Rbbr83 netL83 node_4 -1218.5657470763852
Cbr83 netL83 node_4 -5.720744164010576e-19

* Branch 84
Rabr84 node_2 netRa84 17076.407724338933
Lbr84 netRa84 netL84 -3.448861053776215e-12
Rbbr84 netL84 node_4 -18115.06729750464
Cbr84 netL84 node_4 -1.1147925517218202e-20

* Branch 85
Rabr85 node_2 netRa85 2860.046173329609
Lbr85 netRa85 netL85 -2.4629199543177638e-12
Rbbr85 netL85 node_4 -6602.351344102589
Cbr85 netL85 node_4 -1.3037078966549096e-19

* Branch 86
Rabr86 node_2 netRa86 -3102.1243371203204
Lbr86 netRa86 netL86 2.040297340443206e-12
Rbbr86 netL86 node_4 4457.741068763043
Cbr86 netL86 node_4 1.4749148753116585e-19

* Branch 87
Rabr87 node_2 netRa87 1103.6572184777676
Lbr87 netRa87 netL87 -1.3585402975385944e-12
Rbbr87 netL87 node_4 -4214.7477921096815
Cbr87 netL87 node_4 -2.9183628088175393e-19

* Branch 88
Rabr88 node_2 netRa88 361.4797861419759
Lbr88 netRa88 netL88 4.0601780677053033e-13
Rbbr88 netL88 node_4 -1475.8901776766386
Cbr88 netL88 node_4 7.615708925404057e-19

* Branch 89
Rabr89 node_2 netRa89 6459.643934136225
Lbr89 netRa89 netL89 -2.671616447030169e-12
Rbbr89 netL89 node_4 -8681.702761175156
Cbr89 netL89 node_4 -4.762567948775816e-20

* Branch 90
Rabr90 node_2 netRa90 305236.4323058897
Lbr90 netRa90 netL90 -8.602976740731104e-12
Rbbr90 netL90 node_4 -305557.20793087635
Cbr90 netL90 node_4 -9.223827753209783e-23

* Branch 91
Rabr91 node_2 netRa91 1712.6314846521911
Lbr91 netRa91 netL91 -1.3398528049181944e-12
Rbbr91 netL91 node_4 -3981.714291525994
Cbr91 netL91 node_4 -1.9637161838710213e-19

* Branch 92
Rabr92 node_2 netRa92 447.20075033942777
Lbr92 netRa92 netL92 -7.321218807381488e-13
Rbbr92 netL92 node_4 -2794.4287257866163
Cbr92 netL92 node_4 -5.85095196734083e-19

* Branch 93
Rabr93 node_2 netRa93 364.07389284885517
Lbr93 netRa93 netL93 -6.843695206288304e-13
Rbbr93 netL93 node_4 -3078.4794038836653
Cbr93 netL93 node_4 -6.094490915581987e-19

* Branch 94
Rabr94 node_2 netRa94 270.114250332611
Lbr94 netRa94 netL94 1.537142347544479e-13
Rbbr94 netL94 node_4 -479.7347203110407
Cbr94 netL94 node_4 1.186958462883246e-18

* Branch 95
Rabr95 node_2 netRa95 3060.4662444092996
Lbr95 netRa95 netL95 -1.2538366100289087e-12
Rbbr95 netL95 node_4 -4198.507923264918
Cbr95 netL95 node_4 -9.75209383945954e-20

* Branch 96
Rabr96 node_2 netRa96 11.705318774402134
Lbr96 netRa96 netL96 -1.1628739433697329e-13
Rbbr96 netL96 node_4 -3109.872753093637
Cbr96 netL96 node_4 -3.0502534725804185e-18

* Branch 97
Rabr97 node_2 netRa97 -40.65528186271221
Lbr97 netRa97 netL97 -8.294983330054942e-14
Rbbr97 netL97 node_4 518.1656623694537
Cbr97 netL97 node_4 -4.005095831521046e-18

* Branch 98
Rabr98 node_2 netRa98 226.4449731379838
Lbr98 netRa98 netL98 -7.620953563083529e-14
Rbbr98 netL98 node_4 -312.6957322020706
Cbr98 netL98 node_4 -1.0544090115377733e-18

* Branch 99
Rabr99 node_2 netRa99 86.65392361926847
Lbr99 netRa99 netL99 -4.54587465616041e-14
Rbbr99 netL99 node_4 -150.45760176059534
Cbr99 netL99 node_4 -3.3705584930474447e-18

.ends


* Y'33
.subckt yp33 node_3 0
* Branch 0
Rabr0 node_3 netRa0 -705962.9055143105
Lbr0 netRa0 netL0 7.724842809707413e-11
Rbbr0 netL0 0 733571.8976533264
Cbr0 netL0 0 1.4851763060980175e-22

* Branch 1
Rabr1 node_3 netRa1 -30432.473174496496
Lbr1 netRa1 netL1 1.6901793382716296e-11
Rbbr1 netL1 0 60559.98662623316
Cbr1 netL1 0 8.988996287688979e-21

* Branch 2
Rabr2 node_3 netRa2 -4371.6695990265835
Lbr2 netRa2 netL2 5.911983327542604e-12
Rbbr2 netL2 0 29500.38670700461
Cbr2 netL2 0 4.406243518899249e-20

* Branch 3
Rabr3 node_3 netRa3 20953.432157082425
Lbr3 netRa3 netL3 -6.187713074345231e-12
Rbbr3 netL3 0 -26971.635104748348
Cbr3 netL3 0 -1.0855684084347603e-20

* Branch 4
Rabr4 node_3 netRa4 5062.304042789573
Lbr4 netRa4 netL4 4.741491032168722e-12
Rbbr4 netL4 0 -19887.35325936312
Cbr4 netL4 0 4.8345277950955904e-20

* Branch 5
Rabr5 node_3 netRa5 -12179599.462676687
Lbr5 netRa5 netL5 2.1705435746798125e-10
Rbbr5 netL5 0 12191603.523825865
Cbr5 netL5 0 1.4612271156301791e-24

* Branch 6
Rabr6 node_3 netRa6 -5154.75687091934
Lbr6 netRa6 netL6 -7.0987785793872514e-12
Rbbr6 netL6 0 23816.7810221942
Cbr6 netL6 0 -5.947085836870857e-20

* Branch 7
Rabr7 node_3 netRa7 -1806.3393879868672
Lbr7 netRa7 netL7 -4.609000622309771e-12
Rbbr7 netL7 0 29139.741087386556
Cbr7 netL7 0 -9.197509410268532e-20

* Branch 8
Rabr8 node_3 netRa8 -7609.305761187026
Lbr8 netRa8 netL8 -8.431985130953775e-12
Rbbr8 netL8 0 24125.362595045335
Cbr8 netL8 0 -4.678357770882642e-20

* Branch 9
Rabr9 node_3 netRa9 37199.66484274863
Lbr9 netRa9 netL9 -2.6392984742290688e-11
Rbbr9 netL9 0 -64745.2583870525
Cbr9 netL9 0 -1.083329151732874e-20

* Branch 10
Rabr10 node_3 netRa10 -4949.559155009403
Lbr10 netRa10 netL10 -6.728877294079904e-12
Rbbr10 netL10 0 23387.24799880445
Cbr10 netL10 0 -5.940096247823609e-20

* Branch 11
Rabr11 node_3 netRa11 186.96987715184088
Lbr11 netRa11 netL11 -5.043690907116664e-12
Rbbr11 netL11 0 -217139.9801052822
Cbr11 netL11 0 -8.744149716888656e-20

* Branch 12
Rabr12 node_3 netRa12 -4443.232998128944
Lbr12 netRa12 netL12 -2.346254147666788e-11
Rbbr12 netL12 0 79450.71270918466
Cbr12 netL12 0 -7.169940026578391e-20

* Branch 13
Rabr13 node_3 netRa13 -15683.93100152351
Lbr13 netRa13 netL13 -1.4580551908369822e-11
Rbbr13 netL13 0 36894.644357079225
Cbr13 netL13 0 -2.5516999990492088e-20

* Branch 14
Rabr14 node_3 netRa14 -21076.0651566328
Lbr14 netRa14 netL14 -1.2412641694614614e-11
Rbbr14 netL14 0 33314.312696347275
Cbr14 netL14 0 -1.781944791479807e-20

* Branch 15
Rabr15 node_3 netRa15 -2058.1650580893206
Lbr15 netRa15 netL15 -1.0159017088692977e-11
Rbbr15 netL15 0 58896.73731662614
Cbr15 netL15 0 -8.960413872403252e-20

* Branch 16
Rabr16 node_3 netRa16 744079.0579405786
Lbr16 netRa16 netL16 -6.52450917150985e-11
Rbbr16 netL16 0 -763870.3448830768
Cbr16 netL16 0 -1.146610720044233e-22

* Branch 17
Rabr17 node_3 netRa17 367574.23153761815
Lbr17 netRa17 netL17 -9.968650524032659e-11
Rbbr17 netL17 0 -381588.52924835065
Cbr17 netL17 0 -7.083016810607213e-22

* Branch 18
Rabr18 node_3 netRa18 -2112.673122711461
Lbr18 netRa18 netL18 -1.3481240339407883e-11
Rbbr18 netL18 0 73844.3988448953
Cbr18 netL18 0 -9.390747783849951e-20

* Branch 19
Rabr19 node_3 netRa19 -205952.94232902565
Lbr19 netRa19 netL19 -4.8506791757999134e-11
Rbbr19 netL19 0 239914.42982606613
Cbr19 netL19 0 -9.84480154304695e-22

* Branch 20
Rabr20 node_3 netRa20 12393.053956764776
Lbr20 netRa20 netL20 1.9360943397498247e-11
Rbbr20 netL20 0 -25630.566101896315
Cbr20 netL20 0 6.211193252336146e-20

* Branch 21
Rabr21 node_3 netRa21 2057.044560152808
Lbr21 netRa21 netL21 -1.0104162959112472e-11
Rbbr21 netL21 0 -77405.60028161522
Cbr21 netL21 0 -5.994589821577561e-20

* Branch 22
Rabr22 node_3 netRa22 -11931.618513503283
Lbr22 netRa22 netL22 -1.5515229626272288e-11
Rbbr22 netL22 0 39403.30344736488
Cbr22 netL22 0 -3.349547043787389e-20

* Branch 23
Rabr23 node_3 netRa23 2994.954441656832
Lbr23 netRa23 netL23 -4.898444415819764e-12
Rbbr23 netL23 0 -24510.205672656964
Cbr23 netL23 0 -6.553732012572713e-20

* Branch 24
Rabr24 node_3 netRa24 60075.74470668897
Lbr24 netRa24 netL24 -6.560192344755578e-11
Rbbr24 netL24 0 -88396.4634263515
Cbr24 netL24 0 -1.221159900631969e-20

* Branch 25
Rabr25 node_3 netRa25 -170.3381965672079
Lbr25 netRa25 netL25 -4.361681264999382e-12
Rbbr25 netL25 0 370257.4089953235
Cbr25 netL25 0 -9.40391505929853e-20

* Branch 26
Rabr26 node_3 netRa26 2454.0379322916365
Lbr26 netRa26 netL26 -1.147709490058005e-11
Rbbr26 netL26 0 -73950.01869855393
Cbr26 netL26 0 -6.049554170794187e-20

* Branch 27
Rabr27 node_3 netRa27 106512.33625827209
Lbr27 netRa27 netL27 -4.915566888404193e-11
Rbbr27 netL27 0 -116525.10138766577
Cbr27 netL27 0 -3.9440310181597706e-21

* Branch 28
Rabr28 node_3 netRa28 -682757.047932897
Lbr28 netRa28 netL28 -4.5958425746290715e-11
Rbbr28 netL28 0 691972.7456909094
Cbr28 netL28 0 -9.73360085886382e-23

* Branch 29
Rabr29 node_3 netRa29 -3598.5857088223647
Lbr29 netRa29 netL29 -1.52752070459731e-11
Rbbr29 netL29 0 50500.06162435705
Cbr29 netL29 0 -8.739802604767359e-20

* Branch 30
Rabr30 node_3 netRa30 1105.5831481642936
Lbr30 netRa30 netL30 -1.13526120938536e-11
Rbbr30 netL30 0 -66816.7094803937
Cbr30 netL30 0 -1.410513693117661e-19

* Branch 31
Rabr31 node_3 netRa31 -12886.912629231318
Lbr31 netRa31 netL31 -2.93010076141139e-11
Rbbr31 netL31 0 56239.11690217188
Cbr31 netL31 0 -4.1230783634198917e-20

* Branch 32
Rabr32 node_3 netRa32 192754.6598563173
Lbr32 netRa32 netL32 -5.014249003427237e-11
Rbbr32 netL32 0 -209925.49367011886
Cbr32 netL32 0 -1.2364407703953339e-21

* Branch 33
Rabr33 node_3 netRa33 -9710.062717933359
Lbr33 netRa33 netL33 -1.1891585538731186e-11
Rbbr33 netL33 0 30621.389039119404
Cbr33 netL33 0 -4.039708377990733e-20

* Branch 34
Rabr34 node_3 netRa34 344583.9489549469
Lbr34 netRa34 netL34 -1.0352907114870265e-10
Rbbr34 netL34 0 -384237.4120280446
Cbr34 netL34 0 -7.801899947451745e-22

* Branch 35
Rabr35 node_3 netRa35 -4096.969979014337
Lbr35 netRa35 netL35 -5.818164891527988e-12
Rbbr35 netL35 0 21605.370118112936
Cbr35 netL35 0 -6.638084509385841e-20

* Branch 36
Rabr36 node_3 netRa36 -2581.521967127217
Lbr36 netRa36 netL36 -1.2126246197830055e-11
Rbbr36 netL36 0 55469.87505326275
Cbr36 netL36 0 -8.747651075300893e-20

* Branch 37
Rabr37 node_3 netRa37 12660.211824620268
Lbr37 netRa37 netL37 -9.668188991345223e-12
Rbbr37 netL37 0 -34139.46400298232
Cbr37 netL37 0 -2.2256804210081553e-20

* Branch 38
Rabr38 node_3 netRa38 42723.94625185669
Lbr38 netRa38 netL38 -3.560919958851308e-11
Rbbr38 netL38 0 -57186.52363472678
Cbr38 netL38 0 -1.450234437203997e-20

* Branch 39
Rabr39 node_3 netRa39 -56779.41167204522
Lbr39 netRa39 netL39 -1.430901562969061e-11
Rbbr39 netL39 0 68291.80976265944
Cbr39 netL39 0 -3.6954716414301496e-21

* Branch 40
Rabr40 node_3 netRa40 -10372.490317897114
Lbr40 netRa40 netL40 -3.321045627464354e-11
Rbbr40 netL40 0 64004.40072724727
Cbr40 netL40 0 -5.08993016078426e-20

* Branch 41
Rabr41 node_3 netRa41 -93393.32285811004
Lbr41 netRa41 netL41 3.148263704257914e-11
Rbbr41 netL41 0 117546.41528175879
Cbr41 netL41 0 2.8627455100775782e-21

* Branch 42
Rabr42 node_3 netRa42 -4259.547476559263
Lbr42 netRa42 netL42 -1.3936395820028126e-11
Rbbr42 netL42 0 43802.696878489514
Cbr42 netL42 0 -7.591504349914567e-20

* Branch 43
Rabr43 node_3 netRa43 -875.9634629704551
Lbr43 netRa43 netL43 -3.8474632243090216e-12
Rbbr43 netL43 0 45718.09360847983
Cbr43 netL43 0 -9.809392633506256e-20

* Branch 44
Rabr44 node_3 netRa44 72430580.83444947
Lbr44 netRa44 netL44 -1.4457725195146906e-09
Rbbr44 netL44 0 -72474855.67711994
Cbr44 netL44 0 -2.7540156299254255e-25

* Branch 45
Rabr45 node_3 netRa45 1941224.6398812428
Lbr45 netRa45 netL45 -3.5757469294803664e-10
Rbbr45 netL45 0 -1971938.5130898138
Cbr45 netL45 0 -9.336736327074235e-23

* Branch 46
Rabr46 node_3 netRa46 67837.33835132401
Lbr46 netRa46 netL46 -5.3307297310132544e-11
Rbbr46 netL46 0 -116347.98424490231
Cbr46 netL46 0 -6.741345579929173e-21

* Branch 47
Rabr47 node_3 netRa47 -3505.370860922201
Lbr47 netRa47 netL47 -1.2195731904390581e-11
Rbbr47 netL47 0 44592.09184153942
Cbr47 netL47 0 -7.865023627678333e-20

* Branch 48
Rabr48 node_3 netRa48 532496.3047084453
Lbr48 netRa48 netL48 -2.074283703705041e-10
Rbbr48 netL48 0 -576303.1513319083
Cbr48 netL48 0 -6.754076083820524e-22

* Branch 49
Rabr49 node_3 netRa49 327577.4195008809
Lbr49 netRa49 netL49 1.5325810748630103e-10
Rbbr49 netL49 0 -464949.5109429585
Cbr49 netL49 0 1.0071636848888382e-21

* Branch 50
Rabr50 node_3 netRa50 1158949.329667559
Lbr50 netRa50 netL50 1.9668623534212353e-10
Rbbr50 netL50 0 -1227877.262791389
Cbr50 netL50 0 1.38254436161034e-22

* Branch 51
Rabr51 node_3 netRa51 -6785.627511166113
Lbr51 netRa51 netL51 2.7696917550220495e-10
Rbbr51 netL51 0 18850520.59303113
Cbr51 netL51 0 2.0422973748803988e-21

* Branch 52
Rabr52 node_3 netRa52 -107201.00137912108
Lbr52 netRa52 netL52 3.0029608252007965e-11
Rbbr52 netL52 0 127754.07989070888
Cbr52 netL52 0 2.191797133658209e-21

* Branch 53
Rabr53 node_3 netRa53 -36707997.557124995
Lbr53 netRa53 netL53 -1.0495372867180703e-09
Rbbr53 netL53 0 36778264.24513986
Cbr53 netL53 0 -7.774343691823666e-25

* Branch 54
Rabr54 node_3 netRa54 -273419.6106628902
Lbr54 netRa54 netL54 -1.515291752188925e-10
Rbbr54 netL54 0 497749.77841055754
Cbr54 netL54 0 -1.114257988411585e-21

* Branch 55
Rabr55 node_3 netRa55 -514093.03762860654
Lbr55 netRa55 netL55 -7.399724988806406e-11
Rbbr55 netL55 0 541927.8441979771
Cbr55 netL55 0 -2.6565368806720886e-22

* Branch 56
Rabr56 node_3 netRa56 717719.5289267235
Lbr56 netRa56 netL56 -2.706859877618404e-10
Rbbr56 netL56 0 -800090.7919152303
Cbr56 netL56 0 -4.711478947387428e-22

* Branch 57
Rabr57 node_3 netRa57 3867699.2024979633
Lbr57 netRa57 netL57 -6.75131774920356e-10
Rbbr57 netL57 0 -3955264.6716341916
Cbr57 netL57 0 -4.4123743537326937e-23

* Branch 58
Rabr58 node_3 netRa58 1540673.319843689
Lbr58 netRa58 netL58 6.90792943646239e-10
Rbbr58 netL58 0 -1780818.6657076464
Cbr58 netL58 0 2.5190862493639864e-22

* Branch 59
Rabr59 node_3 netRa59 -502982.30711073795
Lbr59 netRa59 netL59 -4.86898506930169e-11
Rbbr59 netL59 0 515899.5436079717
Cbr59 netL59 0 -1.876577657537604e-22

* Branch 60
Rabr60 node_3 netRa60 117813506.32014336
Lbr60 netRa60 netL60 -3.080293847219002e-09
Rbbr60 netL60 0 -117881107.16001149
Cbr60 netL60 0 -2.217896029298844e-25

* Branch 61
Rabr61 node_3 netRa61 843988.4160438213
Lbr61 netRa61 netL61 -2.9681318568594904e-10
Rbbr61 netL61 0 -961140.6097250925
Cbr61 netL61 0 -3.6577463419359934e-22

* Branch 62
Rabr62 node_3 netRa62 298443.5432245906
Lbr62 netRa62 netL62 -2.45350247724453e-10
Rbbr62 netL62 0 -442156.1573504256
Cbr62 netL62 0 -1.8578465462480703e-21

* Branch 63
Rabr63 node_3 netRa63 1356656.9401296503
Lbr63 netRa63 netL63 -5.008392944695289e-10
Rbbr63 netL63 0 -1461747.6905067447
Cbr63 netL63 0 -2.5246814011775205e-22

* Branch 64
Rabr64 node_3 netRa64 2847711.0395825882
Lbr64 netRa64 netL64 -5.456082014218568e-10
Rbbr64 netL64 0 -2946015.5421454064
Cbr64 netL64 0 -6.502495119570192e-23

* Branch 65
Rabr65 node_3 netRa65 14815917.064358367
Lbr65 netRa65 netL65 1.2928437026017643e-09
Rbbr65 netL65 0 -14994067.150580825
Cbr65 netL65 0 5.820082904937985e-24

* Branch 66
Rabr66 node_3 netRa66 3680229.1410724334
Lbr66 netRa66 netL66 -8.486468143237895e-10
Rbbr66 netL66 0 -3813815.38343749
Cbr66 netL66 0 -6.045197087938148e-23

* Branch 67
Rabr67 node_3 netRa67 -116489.6369226275
Lbr67 netRa67 netL67 1.0233752665032934e-10
Rbbr67 netL67 0 224199.38027541287
Cbr67 netL67 0 3.9157850037986036e-21

* Branch 68
Rabr68 node_3 netRa68 -2227.494749921022
Lbr68 netRa68 netL68 -9.847938799496818e-12
Rbbr68 netL68 0 53668.58111603286
Cbr68 netL68 0 -8.26404168528989e-20

* Branch 69
Rabr69 node_3 netRa69 373933.8931488857
Lbr69 netRa69 netL69 -2.9971702109555133e-10
Rbbr69 netL69 0 -516961.18957320607
Cbr69 netL69 0 -1.5496529721338953e-21

* Branch 70
Rabr70 node_3 netRa70 -20794.327878914162
Lbr70 netRa70 netL70 -2.336391721185464e-10
Rbbr70 netL70 0 2408765.3037501005
Cbr70 netL70 0 -4.6843072441569295e-21

* Branch 71
Rabr71 node_3 netRa71 -289110.1579816158
Lbr71 netRa71 netL71 -5.817888567487418e-11
Rbbr71 netL71 0 318485.54104531783
Cbr71 netL71 0 -6.318936089293876e-22

* Branch 72
Rabr72 node_3 netRa72 296778.2861814873
Lbr72 netRa72 netL72 -2.737440221313413e-10
Rbbr72 netL72 0 -516917.5096068864
Cbr72 netL72 0 -1.783904981319676e-21

* Branch 73
Rabr73 node_3 netRa73 2300738.796462884
Lbr73 netRa73 netL73 1.7370885129143776e-09
Rbbr73 netL73 0 -3579587.1630521226
Cbr73 netL73 0 2.1096284909060346e-22

* Branch 74
Rabr74 node_3 netRa74 -95141.25438792603
Lbr74 netRa74 netL74 -4.795411333043941e-11
Rbbr74 netL74 0 162597.6350757036
Cbr74 netL74 0 -3.1000821471157706e-21

* Branch 75
Rabr75 node_3 netRa75 -850.0775022184781
Lbr75 netRa75 netL75 -9.610285876734209e-12
Rbbr75 netL75 0 130091.31769909587
Cbr75 netL75 0 -8.695042754913689e-20

* Branch 76
Rabr76 node_3 netRa76 -132617447.36328721
Lbr76 netRa76 netL76 7.642124097212954e-09
Rbbr76 netL76 0 133667241.40890834
Cbr76 netL76 0 4.311100425286997e-25

* Branch 77
Rabr77 node_3 netRa77 181310.05695974143
Lbr77 netRa77 netL77 -3.9289333035346267e-10
Rbbr77 netL77 0 -1041545.7451291383
Cbr77 netL77 0 -2.080394367614805e-21

* Branch 78
Rabr78 node_3 netRa78 798124.1683924231
Lbr78 netRa78 netL78 -4.5330166072321707e-10
Rbbr78 netL78 0 -966425.509727555
Cbr78 netL78 0 -5.87667454346288e-22

* Branch 79
Rabr79 node_3 netRa79 -168826.05670789225
Lbr79 netRa79 netL79 7.311608054008849e-10
Rbbr79 netL79 0 3601292.3455465143
Cbr79 netL79 0 1.2020986132683026e-21

* Branch 80
Rabr80 node_3 netRa80 2096165.4432333275
Lbr80 netRa80 netL80 -7.07665779936912e-10
Rbbr80 netL80 0 -2346276.326563179
Cbr80 netL80 0 -1.4388079819563217e-22

* Branch 81
Rabr81 node_3 netRa81 488884.712362349
Lbr81 netRa81 netL81 4.197715432666388e-10
Rbbr81 netL81 0 -1142440.6031623795
Cbr81 netL81 0 7.5169714744596015e-22

* Branch 82
Rabr82 node_3 netRa82 226251.86844363727
Lbr82 netRa82 netL82 2.4667030607325185e-10
Rbbr82 netL82 0 -753706.5416117541
Cbr82 netL82 0 1.4468117299453752e-21

* Branch 83
Rabr83 node_3 netRa83 35950.67836228122
Lbr83 netRa83 netL83 1.441497579538746e-10
Rbbr83 netL83 0 -1029856.5301805594
Cbr83 netL83 0 3.897416103653704e-21

* Branch 84
Rabr84 node_3 netRa84 48852.76307388455
Lbr84 netRa84 netL84 1.5531585589106034e-10
Rbbr84 netL84 0 -969057.6943752544
Cbr84 netL84 0 3.2839880314989384e-21

* Branch 85
Rabr85 node_3 netRa85 160168.67886141955
Lbr85 netRa85 netL85 2.2204384818175008e-10
Rbbr85 netL85 0 -779613.4724914046
Cbr85 netL85 0 1.778974394308643e-21

* Branch 86
Rabr86 node_3 netRa86 -196017.10956789483
Lbr86 netRa86 netL86 9.706714946986738e-11
Rbbr86 netL86 0 318803.8132629148
Cbr86 netL86 0 1.5530561421407492e-21

* Branch 87
Rabr87 node_3 netRa87 57907275.603111885
Lbr87 netRa87 netL87 -3.927005944481687e-09
Rbbr87 netL87 0 -58269932.10705824
Cbr87 netL87 0 -1.163789662671198e-24

* Branch 88
Rabr88 node_3 netRa88 -121766.48419097858
Lbr88 netRa88 netL88 1.4441029655673356e-10
Rbbr88 netL88 0 483826.3043723821
Cbr88 netL88 0 2.4501801952591272e-21

* Branch 89
Rabr89 node_3 netRa89 316866.67816753377
Lbr89 netRa89 netL89 1.843655554688169e-10
Rbbr89 netL89 0 -549375.0921755288
Cbr89 netL89 0 1.0593124168570997e-21

* Branch 90
Rabr90 node_3 netRa90 -276869.22555163916
Lbr90 netRa90 netL90 -5.675059289387417e-11
Rbbr90 netL90 0 310820.8167138067
Cbr90 netL90 0 -6.59505259972059e-22

* Branch 91
Rabr91 node_3 netRa91 -54360.55232602933
Lbr91 netRa91 netL91 5.287316536714747e-11
Rbbr91 netL91 0 140375.30157294575
Cbr91 netL91 0 6.92620994770501e-21

* Branch 92
Rabr92 node_3 netRa92 -93316.35847724618
Lbr92 netRa92 netL92 -3.9424906355186915e-11
Rbbr92 netL92 0 140860.68729870924
Cbr92 netL92 0 -2.9999394916798885e-21

* Branch 93
Rabr93 node_3 netRa93 -2559.8793797866524
Lbr93 netRa93 netL93 -3.8309286709708616e-12
Rbbr93 netL93 0 21217.83131968205
Cbr93 netL93 0 -7.058865399519185e-20

* Branch 94
Rabr94 node_3 netRa94 1583632.1360505063
Lbr94 netRa94 netL94 3.2311644310110723e-10
Rbbr94 netL94 0 -1678906.9371145773
Cbr94 netL94 0 1.2154281895460292e-22

* Branch 95
Rabr95 node_3 netRa95 590039.0473009644
Lbr95 netRa95 netL95 3.8542306057829296e-10
Rbbr95 netL95 0 -901905.6305815689
Cbr95 netL95 0 7.245527833556167e-22

* Branch 96
Rabr96 node_3 netRa96 4024.978381589201
Lbr96 netRa96 netL96 5.9150886999369e-12
Rbbr96 netL96 0 -30143.949140004075
Cbr96 netL96 0 4.8798695231469904e-20

* Branch 97
Rabr97 node_3 netRa97 53110.23937755876
Lbr97 netRa97 netL97 7.261902548753509e-11
Rbbr97 netL97 0 -273781.9946919963
Cbr97 netL97 0 4.999005776901391e-21

* Branch 98
Rabr98 node_3 netRa98 -121524.26241130641
Lbr98 netRa98 netL98 -4.451688707155523e-11
Rbbr98 netL98 0 179172.7131159494
Cbr98 netL98 0 -2.0464968713422133e-21

* Branch 99
Rabr99 node_3 netRa99 -998.6228412993662
Lbr99 netRa99 netL99 2.4759551337065084e-12
Rbbr99 netL99 0 20047.10852263619
Cbr99 netL99 0 1.174009277689423e-19

.ends


* Y'34
.subckt yp34 node_3 node_4
* Branch 0
Rabr0 node_3 netRa0 -26.463022853310555
Lbr0 netRa0 netL0 -1.0037190454069066e-13
Rbbr0 netL0 node_4 656.0938275224627
Cbr0 netL0 node_4 -1.0985948926513763e-17

* Branch 1
Rabr1 node_3 netRa1 -1105.8031063308663
Lbr1 netRa1 netL1 3.2602274491443213e-13
Rbbr1 netL1 node_4 1360.9090562501021
Cbr1 netL1 node_4 2.114698697234861e-19

* Branch 2
Rabr2 node_3 netRa2 -25.104755952527576
Lbr2 netRa2 netL2 -1.0209513338844321e-13
Rbbr2 netL2 node_4 507.6143916381877
Cbr2 netL2 node_4 -1.1117638416472453e-17

* Branch 3
Rabr3 node_3 netRa3 -23.048606167914834
Lbr3 netRa3 netL3 -1.0662821333129508e-13
Rbbr3 netL3 node_4 501.42358744113193
Cbr3 netL3 node_4 -1.2258300285380828e-17

* Branch 4
Rabr4 node_3 netRa4 -26191.580279530495
Lbr4 netRa4 netL4 1.522653621349258e-12
Rbbr4 netL4 node_4 26432.138891202176
Cbr4 netL4 node_4 2.192760344447124e-21

* Branch 5
Rabr5 node_3 netRa5 393.20730229038315
Lbr5 netRa5 netL5 1.3218323976252255e-13
Rbbr5 netL5 node_4 -528.6873374375763
Cbr5 netL5 node_4 6.468388030531386e-19

* Branch 6
Rabr6 node_3 netRa6 -21.17502570579826
Lbr6 netRa6 netL6 -1.0740644861563358e-13
Rbbr6 netL6 node_4 507.75296985422483
Cbr6 netL6 node_4 -1.2737413883579828e-17

* Branch 7
Rabr7 node_3 netRa7 5282.1075436852325
Lbr7 netRa7 netL7 1.0506056928137687e-12
Rbbr7 netL7 node_4 -5863.120550175992
Cbr7 netL7 node_4 3.4177652087573797e-20

* Branch 8
Rabr8 node_3 netRa8 3352.928347038642
Lbr8 netRa8 netL8 -4.726392063126069e-13
Rbbr8 netL8 node_4 -3550.39403801129
Cbr8 netL8 node_4 -3.950101453480832e-20

* Branch 9
Rabr9 node_3 netRa9 -2811.6583696951925
Lbr9 netRa9 netL9 1.3818833451638938e-13
Rbbr9 netL9 node_4 2834.7749369013823
Cbr9 netL9 node_4 1.7307640824600428e-20

* Branch 10
Rabr10 node_3 netRa10 274.43553119073204
Lbr10 netRa10 netL10 -5.755459072194649e-13
Rbbr10 netL10 node_4 -3841.5607420127594
Cbr10 netL10 node_4 -5.092254050436883e-19

* Branch 11
Rabr11 node_3 netRa11 -207.98314243013726
Lbr11 netRa11 netL11 1.6679963302152373e-13
Rbbr11 netL11 node_4 573.76565738389
Cbr11 netL11 node_4 1.3629248331680192e-18

* Branch 12
Rabr12 node_3 netRa12 509.10725077138426
Lbr12 netRa12 netL12 -4.600595900579927e-13
Rbbr12 netL12 node_4 -1829.7767139442744
Cbr12 netL12 node_4 -4.801374072016169e-19

* Branch 13
Rabr13 node_3 netRa13 -192.2811157557132
Lbr13 netRa13 netL13 -3.194877326342125e-13
Rbbr13 netL13 node_4 1911.6822159319663
Cbr13 netL13 node_4 -9.171767271460916e-19

* Branch 14
Rabr14 node_3 netRa14 124.16562401936454
Lbr14 netRa14 netL14 -5.966612699012101e-14
Rbbr14 netL14 node_4 -221.69195251753857
Cbr14 netL14 node_4 -2.1354887822132506e-18

* Branch 15
Rabr15 node_3 netRa15 -22.052181727191453
Lbr15 netRa15 netL15 -1.0799781987401954e-13
Rbbr15 netL15 node_4 470.45324204052633
Cbr15 netL15 node_4 -1.2268021490290029e-17

* Branch 16
Rabr16 node_3 netRa16 -214.9976210333474
Lbr16 netRa16 netL16 6.398052478902865e-14
Rbbr16 netL16 node_4 279.42288320730165
Cbr16 netL16 node_4 1.0553481213343807e-18

* Branch 17
Rabr17 node_3 netRa17 -6210.7038047640945
Lbr17 netRa17 netL17 -7.341969635563051e-13
Rbbr17 netL17 node_4 6465.989207518655
Cbr17 netL17 node_4 -1.8348828289769125e-20

* Branch 18
Rabr18 node_3 netRa18 18.220176979848397
Lbr18 netRa18 netL18 -3.0357890762327636e-14
Rbbr18 netL18 node_4 -183.21610672606442
Cbr18 netL18 node_4 -8.697763927722289e-18

* Branch 19
Rabr19 node_3 netRa19 36.71325297512373
Lbr19 netRa19 netL19 -9.385519913016021e-14
Rbbr19 netL19 node_4 -498.9342064165094
Cbr19 netL19 node_4 -4.816010117087566e-18

* Branch 20
Rabr20 node_3 netRa20 47.13521958352132
Lbr20 netRa20 netL20 1.0757503596435659e-13
Rbbr20 netL20 node_4 -730.0513444607724
Cbr20 netL20 node_4 3.299967511282423e-18

* Branch 21
Rabr21 node_3 netRa21 640.9200526809711
Lbr21 netRa21 netL21 -2.5861682816134334e-13
Rbbr21 netL21 node_4 -877.055529066115
Cbr21 netL21 node_4 -4.558386876710964e-19

* Branch 22
Rabr22 node_3 netRa22 104.78232259211907
Lbr22 netRa22 netL22 -1.2118328189941644e-13
Rbbr22 netL22 node_4 -404.70966712569776
Cbr22 netL22 node_4 -2.7850380729980926e-18

* Branch 23
Rabr23 node_3 netRa23 4755.745423590554
Lbr23 netRa23 netL23 7.468660005538799e-13
Rbbr23 netL23 node_4 -5087.931627003184
Cbr23 netL23 node_4 3.09676609875986e-20

* Branch 24
Rabr24 node_3 netRa24 -114026.92779420537
Lbr24 netRa24 netL24 2.4865330452408935e-12
Rbbr24 netL24 node_4 114167.33812180346
Cbr24 netL24 node_4 1.9092491245499724e-22

* Branch 25
Rabr25 node_3 netRa25 12.399040180437778
Lbr25 netRa25 netL25 -7.971626001443156e-14
Rbbr25 netL25 node_4 -879.0000427239328
Cbr25 netL25 node_4 -6.532233224222977e-18

* Branch 26
Rabr26 node_3 netRa26 -18.22122999633197
Lbr26 netRa26 netL26 -1.0767051015386673e-13
Rbbr26 netL26 node_4 468.1599779923189
Cbr26 netL26 node_4 -1.4106976318757808e-17

* Branch 27
Rabr27 node_3 netRa27 842.7217446947604
Lbr27 netRa27 netL27 2.3326526821703257e-13
Rbbr27 netL27 node_4 -1061.3059470188846
Cbr27 netL27 node_4 2.621027985493338e-19

* Branch 28
Rabr28 node_3 netRa28 -27069.51091199812
Lbr28 netRa28 netL28 1.9393915016263077e-12
Rbbr28 netL28 node_4 27484.98705679803
Cbr28 netL28 node_4 2.603493136675568e-21

* Branch 29
Rabr29 node_3 netRa29 10246.335271867421
Lbr29 netRa29 netL29 1.2968593762682246e-12
Rbbr29 netL29 node_4 -10646.120683709507
Cbr29 netL29 node_4 1.191363198792843e-20

* Branch 30
Rabr30 node_3 netRa30 2.540550309711882
Lbr30 netRa30 netL30 -9.451657453336078e-14
Rbbr30 netL30 node_4 -3593.52665228352
Cbr30 netL30 node_4 -6.407441048841508e-18

* Branch 31
Rabr31 node_3 netRa31 -18.846870480504712
Lbr31 netRa31 netL31 -8.758946120847414e-14
Rbbr31 netL31 node_4 550.4357947605332
Cbr31 netL31 node_4 -9.043478177067107e-18

* Branch 32
Rabr32 node_3 netRa32 -23.421663100852204
Lbr32 netRa32 netL32 -8.873761379612094e-14
Rbbr32 netL32 node_4 492.1607541865342
Cbr32 netL32 node_4 -8.111699677168469e-18

* Branch 33
Rabr33 node_3 netRa33 577.0248952177922
Lbr33 netRa33 netL33 -4.922717862554037e-13
Rbbr33 netL33 node_4 -1686.1077273463727
Cbr33 netL33 node_4 -5.006489066621096e-19

* Branch 34
Rabr34 node_3 netRa34 7.001241945420931
Lbr34 netRa34 netL34 -8.486800355448287e-14
Rbbr34 netL34 node_4 -1607.8649183448656
Cbr34 netL34 node_4 -6.609279880472802e-18

* Branch 35
Rabr35 node_3 netRa35 18740.033731755266
Lbr35 netRa35 netL35 2.21145636356851e-12
Rbbr35 netL35 node_4 -19488.56841026155
Cbr35 netL35 node_4 6.062406463276418e-21

* Branch 36
Rabr36 node_3 netRa36 -17.148375390745255
Lbr36 netRa36 netL36 -1.213120288569681e-13
Rbbr36 netL36 node_4 486.6288263185043
Cbr36 netL36 node_4 -1.564569741024655e-17

* Branch 37
Rabr37 node_3 netRa37 -1.7013335018188638
Lbr37 netRa37 netL37 -8.309845209008213e-14
Rbbr37 netL37 node_4 11403.122794827406
Cbr37 netL37 node_4 -7.873684724328806e-18

* Branch 38
Rabr38 node_3 netRa38 -21.321217932926572
Lbr38 netRa38 netL38 -1.0666525550592982e-13
Rbbr38 netL38 node_4 517.2557860648542
Cbr38 netL38 node_4 -1.0071099877027843e-17

* Branch 39
Rabr39 node_3 netRa39 195.81758194435443
Lbr39 netRa39 netL39 4.782551548462971e-13
Rbbr39 netL39 node_4 -3693.703527986603
Cbr39 netL39 node_4 6.740097694367996e-19

* Branch 40
Rabr40 node_3 netRa40 -20.074179489581354
Lbr40 netRa40 netL40 -8.649001047541766e-14
Rbbr40 netL40 node_4 550.513651556189
Cbr40 netL40 node_4 -8.080920721276348e-18

* Branch 41
Rabr41 node_3 netRa41 -15.598289125434224
Lbr41 netRa41 netL41 -9.653325409702941e-14
Rbbr41 netL41 node_4 634.3246533980454
Cbr41 netL41 node_4 -1.01811618118434e-17

* Branch 42
Rabr42 node_3 netRa42 -471.32219911355287
Lbr42 netRa42 netL42 -5.031993308467729e-13
Rbbr42 netL42 node_4 1849.5371347135597
Cbr42 netL42 node_4 -5.806094906123526e-19

* Branch 43
Rabr43 node_3 netRa43 -162.6998199541055
Lbr43 netRa43 netL43 6.519323279206408e-13
Rbbr43 netL43 node_4 4475.272362253877
Cbr43 netL43 node_4 8.858840953178494e-19

* Branch 44
Rabr44 node_3 netRa44 -84.65449578846342
Lbr44 netRa44 netL44 -3.527628065488515e-13
Rbbr44 netL44 node_4 1684.2514619892763
Cbr44 netL44 node_4 -2.494706314554129e-18

* Branch 45
Rabr45 node_3 netRa45 -160.85059834443288
Lbr45 netRa45 netL45 1.16228686606064e-12
Rbbr45 netL45 node_4 15214.446684040227
Cbr45 netL45 node_4 4.701191244652874e-19

* Branch 46
Rabr46 node_3 netRa46 -105.03007846020752
Lbr46 netRa46 netL46 5.730653196271971e-13
Rbbr46 netL46 node_4 4865.723267602686
Cbr46 netL46 node_4 1.113133031978516e-18

* Branch 47
Rabr47 node_3 netRa47 11551.325833972103
Lbr47 netRa47 netL47 6.884786769557127e-12
Rbbr47 netL47 node_4 -18597.465388535744
Cbr47 netL47 node_4 3.206751395094529e-20

* Branch 48
Rabr48 node_3 netRa48 -352.3892844499923
Lbr48 netRa48 netL48 -6.442413368629526e-13
Rbbr48 netL48 node_4 3037.7704808337758
Cbr48 netL48 node_4 -6.023148735689535e-19

* Branch 49
Rabr49 node_3 netRa49 765.4509976907697
Lbr49 netRa49 netL49 1.7152084135176343e-12
Rbbr49 netL49 node_4 -8300.132953333927
Cbr49 netL49 node_4 2.702283352032056e-19

* Branch 50
Rabr50 node_3 netRa50 -2094.5781007258333
Lbr50 netRa50 netL50 8.617716484503653e-13
Rbbr50 netL50 node_4 2976.464227972351
Cbr50 netL50 node_4 1.3821797884260674e-19

* Branch 51
Rabr51 node_3 netRa51 7061524.604931917
Lbr51 netRa51 netL51 1.0905747871449284e-10
Rbbr51 netL51 node_4 -7064657.218246907
Cbr51 netL51 node_4 2.1860844500357128e-24

* Branch 52
Rabr52 node_3 netRa52 -9600.195499429183
Lbr52 netRa52 netL52 3.4601684103051357e-12
Rbbr52 netL52 node_4 11802.403443635249
Cbr52 netL52 node_4 3.053725957811532e-20

* Branch 53
Rabr53 node_3 netRa53 5889.718483786015
Lbr53 netRa53 netL53 -4.929367417639151e-12
Rbbr53 netL53 node_4 -12031.753585702389
Cbr53 netL53 node_4 -6.95581436684883e-20

* Branch 54
Rabr54 node_3 netRa54 17460.91358796905
Lbr54 netRa54 netL54 6.188694965902188e-12
Rbbr54 netL54 node_4 -21869.598365230595
Cbr54 netL54 node_4 1.6206678390659186e-20

* Branch 55
Rabr55 node_3 netRa55 1466.8993657415192
Lbr55 netRa55 netL55 1.958196760941988e-12
Rbbr55 netL55 node_4 -6988.25503926285
Cbr55 netL55 node_4 1.9104096530588766e-19

* Branch 56
Rabr56 node_3 netRa56 243.50897657001494
Lbr56 netRa56 netL56 -1.6015278762485378e-12
Rbbr56 netL56 node_4 -5127.888620798584
Cbr56 netL56 node_4 -1.2805615022262096e-18

* Branch 57
Rabr57 node_3 netRa57 239.5031263842592
Lbr57 netRa57 netL57 -1.7962484225662493e-12
Rbbr57 netL57 node_4 -6159.750866341847
Cbr57 netL57 node_4 -1.2153357024478967e-18

* Branch 58
Rabr58 node_3 netRa58 501.3940550147735
Lbr58 netRa58 netL58 8.080588749116678e-13
Rbbr58 netL58 node_4 -2326.89995396317
Cbr58 netL58 node_4 6.928907988873698e-19

* Branch 59
Rabr59 node_3 netRa59 261.619256000243
Lbr59 netRa59 netL59 -1.8838312368697748e-12
Rbbr59 netL59 node_4 -5904.188675594924
Cbr59 netL59 node_4 -1.2172520945914647e-18

* Branch 60
Rabr60 node_3 netRa60 70805.94679176791
Lbr60 netRa60 netL60 -1.508709509152808e-11
Rbbr60 netL60 node_4 -73822.47782399833
Cbr60 netL60 node_4 -2.8861602251141668e-21

* Branch 61
Rabr61 node_3 netRa61 1153.9465555444795
Lbr61 netRa61 netL61 -2.7980809917105314e-12
Rbbr61 netL61 node_4 -4819.6774602588375
Cbr61 netL61 node_4 -5.027128365969279e-19

* Branch 62
Rabr62 node_3 netRa62 403.1701449771649
Lbr62 netRa62 netL62 -1.3346020110444894e-12
Rbbr62 netL62 node_4 -2562.7098061832558
Cbr62 netL62 node_4 -1.2903102981832248e-18

* Branch 63
Rabr63 node_3 netRa63 2269.12744332594
Lbr63 netRa63 netL63 -2.274731233189263e-12
Rbbr63 netL63 node_4 -4489.399037707716
Cbr63 netL63 node_4 -2.2322160458657354e-19

* Branch 64
Rabr64 node_3 netRa64 715.9372955590712
Lbr64 netRa64 netL64 -2.0452291629262206e-12
Rbbr64 netL64 node_4 -4028.6132425542883
Cbr64 netL64 node_4 -7.084114975347396e-19

* Branch 65
Rabr65 node_3 netRa65 641.8704392473098
Lbr65 netRa65 netL65 -2.285325467929816e-12
Rbbr65 netL65 node_4 -3844.498646558833
Cbr65 netL65 node_4 -9.248715519539322e-19

* Branch 66
Rabr66 node_3 netRa66 9631.141707360435
Lbr66 netRa66 netL66 -7.0756743667875986e-12
Rbbr66 netL66 node_4 -15452.854279704967
Cbr66 netL66 node_4 -4.752905979609063e-20

* Branch 67
Rabr67 node_3 netRa67 -4260.427347039759
Lbr67 netRa67 netL67 5.175308077792817e-12
Rbbr67 netL67 node_4 14472.8748380687
Cbr67 netL67 node_4 8.389013360337911e-20

* Branch 68
Rabr68 node_3 netRa68 -62337.18294798937
Lbr68 netRa68 netL68 -1.5101219166412856e-11
Rbbr68 netL68 node_4 68118.71671810752
Cbr68 netL68 node_4 -3.556662173976424e-21

* Branch 69
Rabr69 node_3 netRa69 812.3735880087823
Lbr69 netRa69 netL69 -1.6362494981484036e-12
Rbbr69 netL69 node_4 -2771.4780964073657
Cbr69 netL69 node_4 -7.260878349717944e-19

* Branch 70
Rabr70 node_3 netRa70 4732.095241398282
Lbr70 netRa70 netL70 5.359171693776651e-12
Rbbr70 netL70 node_4 -13507.989996884302
Cbr70 netL70 node_4 8.388334179091835e-20

* Branch 71
Rabr71 node_3 netRa71 6745.9668551315735
Lbr71 netRa71 netL71 -3.653954989807446e-12
Rbbr71 netL71 node_4 -8035.484250196699
Cbr71 netL71 node_4 -6.739045441835596e-20

* Branch 72
Rabr72 node_3 netRa72 4224.710962643614
Lbr72 netRa72 netL72 -2.727580261530639e-12
Rbbr72 netL72 node_4 -5757.0106327884705
Cbr72 netL72 node_4 -1.1211130481428103e-19

* Branch 73
Rabr73 node_3 netRa73 3401.0372673918187
Lbr73 netRa73 netL73 -2.3710136985077433e-12
Rbbr73 netL73 node_4 -4526.404580522324
Cbr73 netL73 node_4 -1.5396587463642546e-19

* Branch 74
Rabr74 node_3 netRa74 4010.988710701119
Lbr74 netRa74 netL74 -3.782692143814445e-12
Rbbr74 netL74 node_4 -8143.3790524683545
Cbr74 netL74 node_4 -1.1575602728387344e-19

* Branch 75
Rabr75 node_3 netRa75 992498.205864703
Lbr75 netRa75 netL75 4.412705773013194e-11
Rbbr75 netL75 node_4 -994013.8114566002
Cbr75 netL75 node_4 4.472935397369945e-23

* Branch 76
Rabr76 node_3 netRa76 -8185.0698105456095
Lbr76 netRa76 netL76 -2.5583974681088725e-12
Rbbr76 netL76 node_4 9714.673431506637
Cbr76 netL76 node_4 -3.218018447664726e-20

* Branch 77
Rabr77 node_3 netRa77 14089.721692040359
Lbr77 netRa77 netL77 4.781337223831186e-12
Rbbr77 netL77 node_4 -14924.612361206573
Cbr77 netL77 node_4 2.2741743458257062e-20

* Branch 78
Rabr78 node_3 netRa78 3064.9308477221552
Lbr78 netRa78 netL78 2.5468556500910123e-12
Rbbr78 netL78 node_4 -7648.998901765406
Cbr78 netL78 node_4 1.0868661408245996e-19

* Branch 79
Rabr79 node_3 netRa79 78348.55896782801
Lbr79 netRa79 netL79 -1.2873699648402413e-11
Rbbr79 netL79 node_4 -80050.14878980494
Cbr79 netL79 node_4 -2.052439264492552e-21

* Branch 80
Rabr80 node_3 netRa80 3826.511901068228
Lbr80 netRa80 netL80 -2.2894071949055295e-12
Rbbr80 netL80 node_4 -5467.03974145268
Cbr80 netL80 node_4 -1.0940101477211582e-19

* Branch 81
Rabr81 node_3 netRa81 22547.966183206412
Lbr81 netRa81 netL81 9.83603923769481e-12
Rbbr81 netL81 node_4 -27036.918034405153
Cbr81 netL81 node_4 1.6138608388250825e-20

* Branch 82
Rabr82 node_3 netRa82 929.230263430972
Lbr82 netRa82 netL82 1.0341604378858076e-12
Rbbr82 netL82 node_4 -1969.913112433275
Cbr82 netL82 node_4 5.65348618358831e-19

* Branch 83
Rabr83 node_3 netRa83 2875.6500279651973
Lbr83 netRa83 netL83 -1.972624758702732e-12
Rbbr83 netL83 node_4 -3718.532867572845
Cbr83 netL83 node_4 -1.843955441591781e-19

* Branch 84
Rabr84 node_3 netRa84 557.8930067956586
Lbr84 netRa84 netL84 1.2110641203385311e-12
Rbbr84 netL84 node_4 -3214.612719595936
Cbr84 netL84 node_4 6.762070025189044e-19

* Branch 85
Rabr85 node_3 netRa85 3587.76673369085
Lbr85 netRa85 netL85 2.1776192141338987e-12
Rbbr85 netL85 node_4 -5223.507700263125
Cbr85 netL85 node_4 1.1624514889563102e-19

* Branch 86
Rabr86 node_3 netRa86 1440246.3528468946
Lbr86 netRa86 netL86 -3.881847773253861e-11
Rbbr86 netL86 node_4 -1440990.1802640476
Cbr86 netL86 node_4 -1.8703921329231652e-23

* Branch 87
Rabr87 node_3 netRa87 10612.250671539716
Lbr87 netRa87 netL87 3.7418662819137585e-12
Rbbr87 netL87 node_4 -11590.553642950586
Cbr87 netL87 node_4 3.0428586997555903e-20

* Branch 88
Rabr88 node_3 netRa88 167068.97397951828
Lbr88 netRa88 netL88 -1.7768777730437835e-11
Rbbr88 netL88 node_4 -168650.92865363354
Cbr88 netL88 node_4 -6.305784457201824e-22

* Branch 89
Rabr89 node_3 netRa89 58133.861737370484
Lbr89 netRa89 netL89 -1.133718251999837e-11
Rbbr89 netL89 node_4 -60958.977963303674
Cbr89 netL89 node_4 -3.1987013692188864e-21

* Branch 90
Rabr90 node_3 netRa90 10187313.292325558
Lbr90 netRa90 netL90 -1.0527173352961239e-10
Rbbr90 netL90 node_4 -10188793.586236265
Cbr90 netL90 node_4 -1.0142053158741605e-24

* Branch 91
Rabr91 node_3 netRa91 -20989.133702607294
Lbr91 netRa91 netL91 5.3246298373224405e-12
Rbbr91 netL91 node_4 23775.38576703332
Cbr91 netL91 node_4 1.0667942468866182e-20

* Branch 92
Rabr92 node_3 netRa92 341.225187980489
Lbr92 netRa92 netL92 5.780492019711906e-13
Rbbr92 netL92 node_4 -1401.4548051928655
Cbr92 netL92 node_4 1.2108672098380169e-18

* Branch 93
Rabr93 node_3 netRa93 15639.403009558533
Lbr93 netRa93 netL93 2.993974993321395e-12
Rbbr93 netL93 node_4 -16395.45422306934
Cbr93 netL93 node_4 1.1678578073962143e-20

* Branch 94
Rabr94 node_3 netRa94 -234.3900463126798
Lbr94 netRa94 netL94 8.641162301665057e-13
Rbbr94 netL94 node_4 7270.276998817867
Cbr94 netL94 node_4 5.050650542620537e-19

* Branch 95
Rabr95 node_3 netRa95 -16898.097054934773
Lbr95 netRa95 netL95 3.086743893815675e-12
Rbbr95 netL95 node_4 18240.57871507494
Cbr95 netL95 node_4 1.0010995780079673e-20

* Branch 96
Rabr96 node_3 netRa96 -239.03172991632755
Lbr96 netRa96 netL96 -4.3951953253359394e-13
Rbbr96 netL96 node_4 2131.965664235314
Cbr96 netL96 node_4 -8.658518107057231e-19

* Branch 97
Rabr97 node_3 netRa97 -33765.35437181658
Lbr97 netRa97 netL97 2.9245980442929683e-12
Rbbr97 netL97 node_4 34381.909785146294
Cbr97 netL97 node_4 2.5185844903991558e-21

* Branch 98
Rabr98 node_3 netRa98 162.46153649464756
Lbr98 netRa98 netL98 3.738478071929244e-14
Rbbr98 netL98 node_4 -192.02554246825807
Cbr98 netL98 node_4 1.2054586293606683e-18

* Branch 99
Rabr99 node_3 netRa99 -1351.9735017379212
Lbr99 netRa99 netL99 3.442442855312887e-13
Rbbr99 netL99 node_4 1583.4348875198202
Cbr99 netL99 node_4 1.5619241232686442e-19

.ends


* Y'44
.subckt yp44 node_4 0
* Branch 0
Rabr0 node_4 netRa0 5498044444.019466
Lbr0 netRa0 netL0 -3.8277347863618727e-08
Rbbr0 netL0 0 -5498862423.882704
Cbr0 netL0 0 -1.2658611377875654e-27

* Branch 1
Rabr1 node_4 netRa1 32184150.931112085
Lbr1 netRa1 netL1 5.845272731540839e-09
Rbbr1 netL1 0 -34482229.466520034
Cbr1 netL1 0 5.290775543791194e-24

* Branch 2
Rabr2 node_4 netRa2 88099111.55998538
Lbr2 netRa2 netL2 3.877374705893374e-09
Rbbr2 netL2 0 -88650341.27809018
Cbr2 netL2 0 4.970011887747448e-25

* Branch 3
Rabr3 node_4 netRa3 2280686905.8931475
Lbr3 netRa3 netL3 4.315169261219721e-08
Rbbr3 netL3 0 -2282645144.30224
Cbr3 netL3 0 8.292460394310792e-27

* Branch 4
Rabr4 node_4 netRa4 1913970.0510267562
Lbr4 netRa4 netL4 -1.4630682709323402e-09
Rbbr4 netL4 0 -3908551.5499597588
Cbr4 netL4 0 -1.923374760961921e-22

* Branch 5
Rabr5 node_4 netRa5 122811856.74348532
Lbr5 netRa5 netL5 1.0910488086357997e-08
Rbbr5 netL5 0 -125004583.41709477
Cbr5 netL5 0 7.120212049903597e-25

* Branch 6
Rabr6 node_4 netRa6 5684462.781610876
Lbr6 netRa6 netL6 8.411494284059904e-10
Rbbr6 netL6 0 -6100118.765993961
Cbr6 netL6 0 2.4332208335355495e-23

* Branch 7
Rabr7 node_4 netRa7 4501706.068570638
Lbr7 netRa7 netL7 2.225116099437697e-09
Rbbr7 netL7 0 -6754509.407272841
Cbr7 netL7 0 7.388808368726602e-23

* Branch 8
Rabr8 node_4 netRa8 4291648.22556679
Lbr8 netRa8 netL8 -2.628833670202595e-09
Rbbr8 netL8 0 -6991364.839576556
Cbr8 netL8 0 -8.659326728926718e-23

* Branch 9
Rabr9 node_4 netRa9 720331470.976051
Lbr9 netRa9 netL9 -1.830179275576975e-08
Rbbr9 netL9 0 -721631115.455015
Cbr9 netL9 0 -3.5191384393889283e-26

* Branch 10
Rabr10 node_4 netRa10 2024062252.7212253
Lbr10 netRa10 netL10 -3.4205839935687545e-08
Rbbr10 netL10 0 -2025588474.438551
Cbr10 netL10 0 -8.340409118175879e-27

* Branch 11
Rabr11 node_4 netRa11 11896635.081236111
Lbr11 netRa11 netL11 -6.310590503661859e-09
Rbbr11 netL11 0 -15806072.475955423
Cbr11 netL11 0 -3.3280586486221833e-23

* Branch 12
Rabr12 node_4 netRa12 994457.2340681334
Lbr12 netRa12 netL12 6.414193080142726e-10
Rbbr12 netL12 0 -1803008.0877982073
Cbr12 netL12 0 3.6123757675320395e-22

* Branch 13
Rabr13 node_4 netRa13 6167133.702135338
Lbr13 netRa13 netL13 -3.4677172721837363e-09
Rbbr13 netL13 0 -9248699.740435405
Cbr13 netL13 0 -6.031527516176343e-23

* Branch 14
Rabr14 node_4 netRa14 12362762.460513495
Lbr14 netRa14 netL14 -6.980570447749425e-09
Rbbr14 netL14 0 -16497400.918999052
Cbr14 netL14 0 -3.395440335085078e-23

* Branch 15
Rabr15 node_4 netRa15 3157583140.0772085
Lbr15 netRa15 netL15 -4.7136837768674086e-08
Rbbr15 netL15 0 -3159350789.8357906
Cbr15 netL15 0 -4.72408652206649e-27

* Branch 16
Rabr16 node_4 netRa16 10657375.766725412
Lbr16 netRa16 netL16 -5.482499423241061e-09
Rbbr16 netL16 0 -14333834.438704483
Cbr16 netL16 0 -3.563902325358899e-23

* Branch 17
Rabr17 node_4 netRa17 12370542.122827433
Lbr17 netRa17 netL17 -7.3878806369085985e-09
Rbbr17 netL17 0 -16655667.287239796
Cbr17 netL17 0 -3.5576471248248407e-23

* Branch 18
Rabr18 node_4 netRa18 11796068.070637127
Lbr18 netRa18 netL18 -6.437834110714678e-09
Rbbr18 netL18 0 -15789583.73477852
Cbr18 netL18 0 -3.4349542436958744e-23

* Branch 19
Rabr19 node_4 netRa19 12334784.744657911
Lbr19 netRa19 netL19 -7.861919040347746e-09
Rbbr19 netL19 0 -16755054.377938012
Cbr19 netL19 0 -3.779092765231325e-23

* Branch 20
Rabr20 node_4 netRa20 11631442.893216966
Lbr20 netRa20 netL20 -8.541324842846456e-09
Rbbr20 netL20 0 -16319348.902251324
Cbr20 netL20 0 -4.4669939783687963e-23

* Branch 21
Rabr21 node_4 netRa21 2029391.4703658405
Lbr21 netRa21 netL21 -5.678269573058815e-10
Rbbr21 netL21 0 -2331120.507871491
Cbr21 netL21 0 -1.1970080771800695e-22

* Branch 22
Rabr22 node_4 netRa22 7790662.935722151
Lbr22 netRa22 netL22 -4.2083741798131226e-09
Rbbr22 netL22 0 -11155379.519617772
Cbr22 netL22 0 -4.817240239870579e-23

* Branch 23
Rabr23 node_4 netRa23 9049115.487628566
Lbr23 netRa23 netL23 -9.820258627902466e-09
Rbbr23 netL23 0 -14166198.345348597
Cbr23 netL23 0 -7.585577519113937e-23

* Branch 24
Rabr24 node_4 netRa24 11794589.668442642
Lbr24 netRa24 netL24 -8.150436452611862e-09
Rbbr24 netL24 0 -16355353.959975779
Cbr24 netL24 0 -4.1988473765409106e-23

* Branch 25
Rabr25 node_4 netRa25 10958419.936401585
Lbr25 netRa25 netL25 -8.851552176324053e-09
Rbbr25 netL25 0 -15747783.791148202
Cbr25 netL25 0 -5.095214828862207e-23

* Branch 26
Rabr26 node_4 netRa26 10081957.299590606
Lbr26 netRa26 netL26 -9.111368918307029e-09
Rbbr26 netL26 0 -15011775.320892993
Cbr26 netL26 0 -5.978001666955536e-23

* Branch 27
Rabr27 node_4 netRa27 9310500.154083405
Lbr27 netRa27 netL27 -4.902522555721876e-09
Rbbr27 netL27 0 -12882790.87113346
Cbr27 netL27 0 -4.070694519987949e-23

* Branch 28
Rabr28 node_4 netRa28 82605504.9116227
Lbr28 netRa28 netL28 -5.4735208576175205e-09
Rbbr28 netL28 0 -83671267.4972111
Cbr28 netL28 0 -7.915876672462875e-25

* Branch 29
Rabr29 node_4 netRa29 9729818.403454734
Lbr29 netRa29 netL29 -9.531349638346282e-09
Rbbr29 netL29 0 -14770243.329670079
Cbr29 netL29 0 -6.593627614345283e-23

* Branch 30
Rabr30 node_4 netRa30 12129661.582027195
Lbr30 netRa30 netL30 -8.913200995449105e-10
Rbbr30 netL30 0 -12356391.550514517
Cbr30 netL30 0 -5.945131380575455e-24

* Branch 31
Rabr31 node_4 netRa31 1581234498.6655872
Lbr31 netRa31 netL31 -3.647087133506949e-08
Rbbr31 netL31 0 -1582718345.9979818
Cbr31 netL31 0 -1.4572627020021226e-26

* Branch 32
Rabr32 node_4 netRa32 8558237.38718418
Lbr32 netRa32 netL32 -1.886093473706167e-09
Rbbr32 netL32 0 -9792999.251676116
Cbr32 netL32 0 -2.2502024875930276e-23

* Branch 33
Rabr33 node_4 netRa33 7042824.714962428
Lbr33 netRa33 netL33 -1.841502987006237e-09
Rbbr33 netL33 0 -8502911.661247257
Cbr33 netL33 0 -3.074849692239873e-23

* Branch 34
Rabr34 node_4 netRa34 -1964256.436485153
Lbr34 netRa34 netL34 3.1769914653301274e-09
Rbbr34 netL34 0 12557923.767423138
Cbr34 netL34 0 1.287334809666206e-22

* Branch 35
Rabr35 node_4 netRa35 3808793.688855279
Lbr35 netRa35 netL35 -1.2340105793997552e-09
Rbbr35 netL35 0 -5046304.576979657
Cbr35 netL35 0 -6.419752710139566e-23

* Branch 36
Rabr36 node_4 netRa36 854318.7174359931
Lbr36 netRa36 netL36 -4.585100761293991e-10
Rbbr36 netL36 0 -1663446.5414106587
Cbr36 netL36 0 -3.22601672942685e-22

* Branch 37
Rabr37 node_4 netRa37 2422456.0078758034
Lbr37 netRa37 netL37 -9.379539697213451e-10
Rbbr37 netL37 0 -3569667.901942922
Cbr37 netL37 0 -1.0845894065881462e-22

* Branch 38
Rabr38 node_4 netRa38 3289649.067140331
Lbr38 netRa38 netL38 -2.6686784089655297e-09
Rbbr38 netL38 0 -6515925.337939366
Cbr38 netL38 0 -1.2448199366057211e-22

* Branch 39
Rabr39 node_4 netRa39 1247310.3280770078
Lbr39 netRa39 netL39 -6.350955809703984e-10
Rbbr39 netL39 0 -2289564.32411752
Cbr39 netL39 0 -2.22368732194194e-22

* Branch 40
Rabr40 node_4 netRa40 7389142.295287981
Lbr40 netRa40 netL40 -8.572075934603152e-09
Rbbr40 netL40 0 -12263116.457037522
Cbr40 netL40 0 -9.458463680929728e-23

* Branch 41
Rabr41 node_4 netRa41 6451373.567151161
Lbr41 netRa41 netL41 -8.460018729804666e-09
Rbbr41 netL41 0 -11613473.144682756
Cbr41 netL41 0 -1.1289645591545212e-22

* Branch 42
Rabr42 node_4 netRa42 4143525.7270509666
Lbr42 netRa42 netL42 -3.4771949974235375e-09
Rbbr42 netL42 0 -7876202.32351917
Cbr42 netL42 0 -1.0653536248771238e-22

* Branch 43
Rabr43 node_4 netRa43 2450250.316101936
Lbr43 netRa43 netL43 -2.3670173664845035e-09
Rbbr43 netL43 0 -6164976.103999941
Cbr43 netL43 0 -1.5668034199399333e-22

* Branch 44
Rabr44 node_4 netRa44 211863.0205791325
Lbr44 netRa44 netL44 -5.841369562460671e-10
Rbbr44 netL44 0 -3209499.9274972375
Cbr44 netL44 0 -8.588523434446736e-22

* Branch 45
Rabr45 node_4 netRa45 2458251.5923600043
Lbr45 netRa45 netL45 -2.471747139239409e-09
Rbbr45 netL45 0 -6271811.61878115
Cbr45 netL45 0 -1.603058627592489e-22

* Branch 46
Rabr46 node_4 netRa46 3102697.2561368784
Lbr46 netRa46 netL46 -6.665903731764887e-09
Rbbr46 netL46 0 -9083504.804443741
Cbr46 netL46 0 -2.364782571170516e-22

* Branch 47
Rabr47 node_4 netRa47 2772751.63795793
Lbr47 netRa47 netL47 -6.0656438535375075e-09
Rbbr47 netL47 0 -8626588.47956454
Cbr47 netL47 0 -2.5354569082662393e-22

* Branch 48
Rabr48 node_4 netRa48 5456614.124029855
Lbr48 netRa48 netL48 -4.846846626075167e-09
Rbbr48 netL48 0 -11499954.02914191
Cbr48 netL48 0 -7.723458092758223e-23

* Branch 49
Rabr49 node_4 netRa49 2579255.008780455
Lbr49 netRa49 netL49 -2.872130454462946e-09
Rbbr49 netL49 0 -6801468.7494954
Cbr49 netL49 0 -1.6371015394260814e-22

* Branch 50
Rabr50 node_4 netRa50 3278763.462294032
Lbr50 netRa50 netL50 -5.678215096238932e-09
Rbbr50 netL50 0 -9413987.342128394
Cbr50 netL50 0 -1.8394229358646038e-22

* Branch 51
Rabr51 node_4 netRa51 6247980.381907658
Lbr51 netRa51 netL51 -2.5687641728994474e-09
Rbbr51 netL51 0 -8708109.564884135
Cbr51 netL51 0 -4.7211709138099936e-23

* Branch 52
Rabr52 node_4 netRa52 2003459.727462485
Lbr52 netRa52 netL52 -2.2928827964160002e-09
Rbbr52 netL52 0 -6147533.93066073
Cbr52 netL52 0 -1.8615322726145445e-22

* Branch 53
Rabr53 node_4 netRa53 2549644.5787758515
Lbr53 netRa53 netL53 -5.095894543519959e-09
Rbbr53 netL53 0 -8618789.29473005
Cbr53 netL53 0 -2.3187146012702746e-22

* Branch 54
Rabr54 node_4 netRa54 4626795.295653279
Lbr54 netRa54 netL54 -1.831575040830936e-09
Rbbr54 netL54 0 -6691665.619041011
Cbr54 netL54 0 -5.915634039309231e-23

* Branch 55
Rabr55 node_4 netRa55 2877495.1684544715
Lbr55 netRa55 netL55 -6.2758798457197944e-09
Rbbr55 netL55 0 -9935056.271921098
Cbr55 netL55 0 -2.195049653921504e-22

* Branch 56
Rabr56 node_4 netRa56 4582867.084529048
Lbr56 netRa56 netL56 -8.761392175403913e-09
Rbbr56 netL56 0 -13655906.217298178
Cbr56 netL56 0 -1.399832508660005e-22

* Branch 57
Rabr57 node_4 netRa57 4527828.442947793
Lbr57 netRa57 netL57 -1.9597095014430045e-09
Rbbr57 netL57 0 -6892238.3780423235
Cbr57 netL57 0 -6.279609910010801e-23

* Branch 58
Rabr58 node_4 netRa58 3121018.6296185986
Lbr58 netRa58 netL58 -3.773357080327225e-09
Rbbr58 netL58 0 -8591874.556891197
Cbr58 netL58 0 -1.407087087403657e-22

* Branch 59
Rabr59 node_4 netRa59 7917646.964567384
Lbr59 netRa59 netL59 -3.048668356295578e-09
Rbbr59 netL59 0 -10847651.334934594
Cbr59 netL59 0 -3.5495326841753546e-23

* Branch 60
Rabr60 node_4 netRa60 1495659.1792975757
Lbr60 netRa60 netL60 -1.874294965205888e-09
Rbbr60 netL60 0 -5419953.339551492
Cbr60 netL60 0 -2.3119934530200477e-22

* Branch 61
Rabr61 node_4 netRa61 2646256.9403818944
Lbr61 netRa61 netL61 -7.673688726209416e-09
Rbbr61 netL61 0 -11430030.034101084
Cbr61 netL61 0 -2.5367502734582076e-22

* Branch 62
Rabr62 node_4 netRa62 2437811.5845753066
Lbr62 netRa62 netL62 -2.8612355685000397e-09
Rbbr62 netL62 0 -7296327.272096502
Cbr62 netL62 0 -1.608534844054799e-22

* Branch 63
Rabr63 node_4 netRa63 2852427.450281576
Lbr63 netRa63 netL63 -3.5074994828542763e-09
Rbbr63 netL63 0 -8195735.506334918
Cbr63 netL63 0 -1.5002926799540463e-22

* Branch 64
Rabr64 node_4 netRa64 441073.5620057562
Lbr64 netRa64 netL64 -1.013666692248911e-09
Rbbr64 netL64 0 -4664262.824761004
Cbr64 netL64 0 -4.926812377637008e-22

* Branch 65
Rabr65 node_4 netRa65 7743894.1913230745
Lbr65 netRa65 netL65 -3.0190900201829792e-09
Rbbr65 netL65 0 -10748820.44448179
Cbr65 netL65 0 -3.627033456248944e-23

* Branch 66
Rabr66 node_4 netRa66 2552106.2729915134
Lbr66 netRa66 netL66 -3.6467070235577275e-09
Rbbr66 netL66 0 -8201725.677091462
Cbr66 netL66 0 -1.7421343819593797e-22

* Branch 67
Rabr67 node_4 netRa67 2956499.679169459
Lbr67 netRa67 netL67 -6.346036473768481e-09
Rbbr67 netL67 0 -11845716.95636326
Cbr67 netL67 0 -1.811940595794971e-22

* Branch 68
Rabr68 node_4 netRa68 1174969.5848849264
Lbr68 netRa68 netL68 -1.6238827686551653e-09
Rbbr68 netL68 0 -5029626.110849511
Cbr68 netL68 0 -2.7477829411895006e-22

* Branch 69
Rabr69 node_4 netRa69 12892980.090991136
Lbr69 netRa69 netL69 -4.526483477104105e-09
Rbbr69 netL69 0 -16681085.034873769
Cbr69 netL69 0 -2.1046545911858504e-23

* Branch 70
Rabr70 node_4 netRa70 2424065.6954499334
Lbr70 netRa70 netL70 -3.943749138685188e-09
Rbbr70 netL70 0 -9142666.542582396
Cbr70 netL70 0 -1.7794494096981316e-22

* Branch 71
Rabr71 node_4 netRa71 2253006.9432776384
Lbr71 netRa71 netL71 -3.878325089772366e-09
Rbbr71 netL71 0 -8762047.321161577
Cbr71 netL71 0 -1.9645807345922508e-22

* Branch 72
Rabr72 node_4 netRa72 2496952.8231511815
Lbr72 netRa72 netL72 -5.930262203934031e-09
Rbbr72 netL72 0 -12101481.745620545
Cbr72 netL72 0 -1.962532156804763e-22

* Branch 73
Rabr73 node_4 netRa73 1294702.9845289888
Lbr73 netRa73 netL73 -3.4465427977347006e-09
Rbbr73 netL73 0 -6512354.4033178715
Cbr73 netL73 0 -4.0875991127225397e-22

* Branch 74
Rabr74 node_4 netRa74 2367596.3741336903
Lbr74 netRa74 netL74 -3.918031520782995e-09
Rbbr74 netL74 0 -8920976.8215822
Cbr74 netL74 0 -1.8549977559380095e-22

* Branch 75
Rabr75 node_4 netRa75 2859855.9204147533
Lbr75 netRa75 netL75 -4.571320573326981e-09
Rbbr75 netL75 0 -11337416.02951457
Cbr75 netL75 0 -1.4098775917023915e-22

* Branch 76
Rabr76 node_4 netRa76 2743466.990077228
Lbr76 netRa76 netL76 -5.6185138752121775e-09
Rbbr76 netL76 0 -12388695.51475675
Cbr76 netL76 0 -1.6530838784700206e-22

* Branch 77
Rabr77 node_4 netRa77 16556813.447232496
Lbr77 netRa77 netL77 -5.926676111417718e-09
Rbbr77 netL77 0 -22094794.351338353
Cbr77 netL77 0 -1.62010766178803e-23

* Branch 78
Rabr78 node_4 netRa78 4568712.08511071
Lbr78 netRa78 netL78 -6.819334657702678e-09
Rbbr78 netL78 0 -12769442.558266435
Cbr78 netL78 0 -1.168888503337303e-22

* Branch 79
Rabr79 node_4 netRa79 3101937.8819239503
Lbr79 netRa79 netL79 -3.936980842147289e-09
Rbbr79 netL79 0 -13930588.507385204
Cbr79 netL79 0 -9.110817903556446e-23

* Branch 80
Rabr80 node_4 netRa80 9511703.648284264
Lbr80 netRa80 netL80 -7.529512677892267e-09
Rbbr80 netL80 0 -14705907.54924851
Cbr80 netL80 0 -5.382876092009291e-23

* Branch 81
Rabr81 node_4 netRa81 4099558.6633277824
Lbr81 netRa81 netL81 -2.5258201459253186e-09
Rbbr81 netL81 0 -7896041.054982219
Cbr81 netL81 0 -7.802861157456962e-23

* Branch 82
Rabr82 node_4 netRa82 4483305.735845635
Lbr82 netRa82 netL82 -3.731962232303364e-09
Rbbr82 netL82 0 -11380792.183607731
Cbr82 netL82 0 -7.314144497304743e-23

* Branch 83
Rabr83 node_4 netRa83 2003704.3164940865
Lbr83 netRa83 netL83 -4.166852508288536e-09
Rbbr83 netL83 0 -20326776.753926482
Cbr83 netL83 0 -1.0230422690372357e-22

* Branch 84
Rabr84 node_4 netRa84 882884870.003833
Lbr84 netRa84 netL84 -6.295258581208615e-08
Rbbr84 netL84 0 -886948510.8017862
Cbr84 netL84 0 -8.039159233500347e-26

* Branch 85
Rabr85 node_4 netRa85 307830338.2519354
Lbr85 netRa85 netL85 -4.467959014875801e-08
Rbbr85 netL85 0 -312447043.2907292
Cbr85 netL85 0 -4.64536468873317e-25

* Branch 86
Rabr86 node_4 netRa86 -5109416.374596926
Lbr86 netRa86 netL86 -3.4862547850938678e-09
Rbbr86 netL86 0 9894175.493700389
Cbr86 netL86 0 -6.896306830049993e-23

* Branch 87
Rabr87 node_4 netRa87 361346586.4920853
Lbr87 netRa87 netL87 3.7892012765364396e-08
Rbbr87 netL87 0 -365804279.6820065
Cbr87 netL87 0 2.86666198416135e-25

* Branch 88
Rabr88 node_4 netRa88 -11703584.290710583
Lbr88 netRa88 netL88 -5.358885413568338e-09
Rbbr88 netL88 0 15045031.783984782
Cbr88 netL88 0 -3.043482581891773e-23

* Branch 89
Rabr89 node_4 netRa89 1093560.9865752084
Lbr89 netRa89 netL89 -7.942320403930404e-10
Rbbr89 netL89 0 -2772315.084328298
Cbr89 netL89 0 -2.6196801006717613e-22

* Branch 90
Rabr90 node_4 netRa90 -11859201.609976321
Lbr90 netRa90 netL90 -2.828769298882514e-09
Rbbr90 netL90 0 13182245.430357434
Cbr90 netL90 0 -1.809497029679172e-23

* Branch 91
Rabr91 node_4 netRa91 13243223.015822481
Lbr91 netRa91 netL91 4.112513906054522e-09
Rbbr91 netL91 0 -16651563.456129402
Cbr91 netL91 0 1.8649443713270384e-23

* Branch 92
Rabr92 node_4 netRa92 6652173.027337104
Lbr92 netRa92 netL92 8.198773961900756e-09
Rbbr92 netL92 0 -14471932.654902054
Cbr92 netL92 0 8.517046085086078e-23

* Branch 93
Rabr93 node_4 netRa93 1443847.1876393394
Lbr93 netRa93 netL93 6.403896519999676e-09
Rbbr93 netL93 0 -22540789.035495006
Cbr93 netL93 0 1.9682407402306576e-22

* Branch 94
Rabr94 node_4 netRa94 -325015.51865675376
Lbr94 netRa94 netL94 4.78917588014708e-09
Rbbr94 netL94 0 66578651.491515405
Cbr94 netL94 0 2.210935434059872e-22

* Branch 95
Rabr95 node_4 netRa95 -27189592.926953506
Lbr95 netRa95 netL95 9.353682256611014e-09
Rbbr95 netL95 0 34507230.80840422
Cbr95 netL95 0 9.96904986519153e-24

* Branch 96
Rabr96 node_4 netRa96 -121979374.89747089
Lbr96 netRa96 netL96 -9.96909023757299e-09
Rbbr96 netL96 0 124202602.28379647
Cbr96 netL96 0 -6.5803395240193305e-25

* Branch 97
Rabr97 node_4 netRa97 176660.09245986477
Lbr97 netRa97 netL97 -7.032667223098798e-11
Rbbr97 netL97 0 -274443.3467020595
Cbr97 netL97 0 -1.4502491898639429e-21

* Branch 98
Rabr98 node_4 netRa98 -278043.8321281024
Lbr98 netRa98 netL98 -2.198303554023032e-10
Rbbr98 netL98 0 862052.0991208036
Cbr98 netL98 0 -9.178315179696557e-22

* Branch 99
Rabr99 node_4 netRa99 -2040307.401834045
Lbr99 netRa99 netL99 4.5579609272628196e-10
Rbbr99 netL99 0 2388619.2275240473
Cbr99 netL99 0 9.348919044865184e-23

.ends


.end
