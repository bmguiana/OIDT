* netlist generated with vector fitting poles and residues

.subckt total_network node_1 node_2 node_3 node_4 
X_11 node_1 0 yp11
X_12 node_1 node_2 yp12
X_13 node_1 node_3 yp13
X_14 node_1 node_4 yp14
X_22 node_2 0 yp22
X_23 node_2 node_3 yp23
X_24 node_2 node_4 yp24
X_33 node_3 0 yp33
X_34 node_3 node_4 yp34
X_44 node_4 0 yp44
.ends


* Y'11
.subckt yp11 node_1 0
* Branch 0
Rabr0 node_1 netRa0 -17434.741458216307
Lbr0 netRa0 netL0 6.740526373739723e-12
Rbbr0 netL0 0 26099.074994125083
Cbr0 netL0 0 1.4549417833506357e-20

* Branch 1
Rabr1 node_1 netRa1 -13712.658527192589
Lbr1 netRa1 netL1 9.591609417966727e-12
Rbbr1 netL1 0 35754.999325864905
Cbr1 netL1 0 1.894519395738335e-20

* Branch 2
Rabr2 node_1 netRa2 144478.16548934887
Lbr2 netRa2 netL2 -2.6722466757353968e-11
Rbbr2 netL2 0 -161146.41183553886
Cbr2 netL2 0 -1.1386218842461405e-21

* Branch 3
Rabr3 node_1 netRa3 8459.185580103274
Lbr3 netRa3 netL3 2.769773287591538e-12
Rbbr3 netL3 0 -11500.42843078262
Cbr3 netL3 0 2.8744330481230347e-20

* Branch 4
Rabr4 node_1 netRa4 58245.77380389142
Lbr4 netRa4 netL4 -3.646357747642789e-11
Rbbr4 netL4 0 -137266.79288243866
Cbr4 netL4 0 -4.490896676445637e-21

* Branch 5
Rabr5 node_1 netRa5 -30655.805703995622
Lbr5 netRa5 netL5 8.873371956305642e-12
Rbbr5 netL5 0 36510.36364210955
Cbr5 netL5 0 7.879355975893072e-21

* Branch 6
Rabr6 node_1 netRa6 -6064.66989393974
Lbr6 netRa6 netL6 6.533446455634442e-12
Rbbr6 netL6 0 19758.641610002323
Cbr6 netL6 0 5.344360400523019e-20

* Branch 7
Rabr7 node_1 netRa7 -11816.268582430588
Lbr7 netRa7 netL7 8.14846499252976e-12
Rbbr7 netL7 0 21433.998439934057
Cbr7 netL7 0 3.1797068402292764e-20

* Branch 8
Rabr8 node_1 netRa8 -23919.82722802769
Lbr8 netRa8 netL8 -1.0150429402726049e-11
Rbbr8 netL8 0 35136.22845276498
Cbr8 netL8 0 -1.216349531338044e-20

* Branch 9
Rabr9 node_1 netRa9 -3205.3186805798073
Lbr9 netRa9 netL9 3.461217409150293e-12
Rbbr9 netL9 0 12953.239912678846
Cbr9 netL9 0 8.190438999478165e-20

* Branch 10
Rabr10 node_1 netRa10 -8025.806705638787
Lbr10 netRa10 netL10 7.988146692544696e-12
Rbbr10 netL10 0 20763.915611366658
Cbr10 netL10 0 4.7165741489186385e-20

* Branch 11
Rabr11 node_1 netRa11 -2428.7784979727626
Lbr11 netRa11 netL11 1.0411366253988582e-11
Rbbr11 netL11 0 51465.60484167352
Cbr11 netL11 0 7.800027492518306e-20

* Branch 12
Rabr12 node_1 netRa12 -64912.90918024948
Lbr12 netRa12 netL12 1.1454909885363925e-11
Rbbr12 netL12 0 70441.81933975346
Cbr12 netL12 0 2.4987869048247227e-21

* Branch 13
Rabr13 node_1 netRa13 107768.13400103145
Lbr13 netRa13 netL13 -4.8916188814723144e-11
Rbbr13 netL13 0 -150073.56390383153
Cbr13 netL13 0 -3.005132874499613e-21

* Branch 14
Rabr14 node_1 netRa14 1494.329860686832
Lbr14 netRa14 netL14 4.160305548389031e-12
Rbbr14 netL14 0 -36081.01434058917
Cbr14 netL14 0 8.034135974950943e-20

* Branch 15
Rabr15 node_1 netRa15 4292.839848094218
Lbr15 netRa15 netL15 -2.5882284250446662e-11
Rbbr15 netL15 0 -167030.33906295954
Cbr15 netL15 0 -3.336296276770568e-20

* Branch 16
Rabr16 node_1 netRa16 -7151.047274606847
Lbr16 netRa16 netL16 -3.3315816896717247e-12
Rbbr16 netL16 0 12181.508133887708
Cbr16 netL16 0 -3.8481454584985896e-20

* Branch 17
Rabr17 node_1 netRa17 -3115.2557725847882
Lbr17 netRa17 netL17 9.958059318132057e-12
Rbbr17 netL17 0 24589.10573980973
Cbr17 netL17 0 1.2478941040161827e-19

* Branch 18
Rabr18 node_1 netRa18 -7321.957269672947
Lbr18 netRa18 netL18 1.073981090872363e-11
Rbbr18 netL18 0 18955.03692131008
Cbr18 netL18 0 7.597448818752743e-20

* Branch 19
Rabr19 node_1 netRa19 -26561.749292795197
Lbr19 netRa19 netL19 1.0303856419627129e-11
Rbbr19 netL19 0 33875.93572525164
Cbr19 netL19 0 1.1397067764686126e-20

* Branch 20
Rabr20 node_1 netRa20 -2909.7167501678955
Lbr20 netRa20 netL20 1.1413144342668333e-11
Rbbr20 netL20 0 42723.773185624996
Cbr20 netL20 0 8.761369663156509e-20

* Branch 21
Rabr21 node_1 netRa21 -662910.2667570976
Lbr21 netRa21 netL21 -3.883175858395346e-11
Rbbr21 netL21 0 668446.8204335788
Cbr21 netL21 0 -8.76951027662842e-23

* Branch 22
Rabr22 node_1 netRa22 6757.307923396253
Lbr22 netRa22 netL22 2.929793441330839e-11
Rbbr22 netL22 0 -120343.87040894774
Cbr22 netL22 0 3.798460875021512e-20

* Branch 23
Rabr23 node_1 netRa23 -9741.997295187613
Lbr23 netRa23 netL23 6.377520699852608e-12
Rbbr23 netL23 0 18370.625444613477
Cbr23 netL23 0 3.536806357454579e-20

* Branch 24
Rabr24 node_1 netRa24 -5025.069348076812
Lbr24 netRa24 netL24 1.2573637012275823e-11
Rbbr24 netL24 0 22088.996242199228
Cbr24 netL24 0 1.1012853653507068e-19

* Branch 25
Rabr25 node_1 netRa25 -8968.615439263032
Lbr25 netRa25 netL25 9.097178175383637e-12
Rbbr25 netL25 0 21961.69985581605
Cbr25 netL25 0 4.5667238972552355e-20

* Branch 26
Rabr26 node_1 netRa26 6903.840246992069
Lbr26 netRa26 netL26 1.2280473393079975e-11
Rbbr26 netL26 0 -62725.7256101052
Cbr26 netL26 0 2.892010637077594e-20

* Branch 27
Rabr27 node_1 netRa27 -11992.441501298865
Lbr27 netRa27 netL27 9.406136025925023e-12
Rbbr27 netL27 0 23157.64423570252
Cbr27 netL27 0 3.358257856640988e-20

* Branch 28
Rabr28 node_1 netRa28 -7497.355604160065
Lbr28 netRa28 netL28 1.2333238513027663e-11
Rbbr28 netL28 0 19682.30495858405
Cbr28 netL28 0 8.214185284800042e-20

* Branch 29
Rabr29 node_1 netRa29 -25172.82463813807
Lbr29 netRa29 netL29 5.359458280322089e-12
Rbbr29 netL29 0 28731.374202973584
Cbr29 netL29 0 7.393513215274594e-21

* Branch 30
Rabr30 node_1 netRa30 3491258.879069282
Lbr30 netRa30 netL30 -1.4224403756691887e-10
Rbbr30 netL30 0 -3508443.848678373
Cbr30 netL30 0 -1.1607965194839369e-23

* Branch 31
Rabr31 node_1 netRa31 -13592.107979259337
Lbr31 netRa31 netL31 6.883402358902737e-12
Rbbr31 netL31 0 21182.929604279994
Cbr31 netL31 0 2.3789127226640474e-20

* Branch 32
Rabr32 node_1 netRa32 -142015.2550429507
Lbr32 netRa32 netL32 3.984186423675544e-11
Rbbr32 netL32 0 147406.1735769769
Cbr32 netL32 0 1.8986143039451915e-21

* Branch 33
Rabr33 node_1 netRa33 -25243.131889176675
Lbr33 netRa33 netL33 1.5000654978998585e-11
Rbbr33 netL33 0 32443.603888339858
Cbr33 netL33 0 1.8228504248035584e-20

* Branch 34
Rabr34 node_1 netRa34 -136456.34560348094
Lbr34 netRa34 netL34 -4.50491874274081e-11
Rbbr34 netL34 0 146523.07104384317
Cbr34 netL34 0 -2.258666230380894e-21

* Branch 35
Rabr35 node_1 netRa35 -4749.448609238146
Lbr35 netRa35 netL35 8.803785387239355e-12
Rbbr35 netL35 0 24727.673302002033
Cbr35 netL35 0 7.395597526004309e-20

* Branch 36
Rabr36 node_1 netRa36 70289.24254578493
Lbr36 netRa36 netL36 -6.984563279240345e-11
Rbbr36 netL36 0 -130859.39707700502
Cbr36 netL36 0 -7.539500845372043e-21

* Branch 37
Rabr37 node_1 netRa37 -26073.446901520212
Lbr37 netRa37 netL37 -6.674887314061092e-12
Rbbr37 netL37 0 31628.27107690573
Cbr37 netL37 0 -8.106938483764605e-21

* Branch 38
Rabr38 node_1 netRa38 -10105.094161469418
Lbr38 netRa38 netL38 1.0472023289747627e-11
Rbbr38 netL38 0 21507.34176402044
Cbr38 netL38 0 4.7884574711969606e-20

* Branch 39
Rabr39 node_1 netRa39 -1645.9652501767148
Lbr39 netRa39 netL39 1.2870166583199347e-11
Rbbr39 netL39 0 49955.20045567157
Cbr39 netL39 0 1.49728370249461e-19

* Branch 40
Rabr40 node_1 netRa40 -8292.491281330413
Lbr40 netRa40 netL40 8.962246367682136e-12
Rbbr40 netL40 0 21239.06319037788
Cbr40 netL40 0 5.058058576639719e-20

* Branch 41
Rabr41 node_1 netRa41 -6069.055567759307
Lbr41 netRa41 netL41 9.849672650715461e-12
Rbbr41 netL41 0 21962.17490450961
Cbr41 netL41 0 7.323759689151003e-20

* Branch 42
Rabr42 node_1 netRa42 35249.47673525623
Lbr42 netRa42 netL42 -6.566371343432593e-11
Rbbr42 netL42 0 -226778.0552024069
Cbr42 netL42 0 -8.140902182860913e-21

* Branch 43
Rabr43 node_1 netRa43 2644.15255505918
Lbr43 netRa43 netL43 1.0925789092444004e-11
Rbbr43 netL43 0 -131086.71635893194
Cbr43 netL43 0 3.2114449314130766e-20

* Branch 44
Rabr44 node_1 netRa44 121444.85688976741
Lbr44 netRa44 netL44 -4.717667711169872e-11
Rbbr44 netL44 0 -176976.51404714314
Cbr44 netL44 0 -2.1917107160755303e-21

* Branch 45
Rabr45 node_1 netRa45 -40854.88172603963
Lbr45 netRa45 netL45 -4.780461387554052e-11
Rbbr45 netL45 0 91741.53923766602
Cbr45 netL45 0 -1.2811175570650372e-20

* Branch 46
Rabr46 node_1 netRa46 99369.92590901478
Lbr46 netRa46 netL46 -8.548309783875094e-11
Rbbr46 netL46 0 -137402.60221627643
Cbr46 netL46 0 -6.241921618761561e-21

* Branch 47
Rabr47 node_1 netRa47 -4356.6866937956165
Lbr47 netRa47 netL47 1.541898849824969e-11
Rbbr47 netL47 0 137070.88269634542
Cbr47 netL47 0 2.5698385314244617e-20

* Branch 48
Rabr48 node_1 netRa48 -83437.7901513481
Lbr48 netRa48 netL48 -1.2520792127573384e-10
Rbbr48 netL48 0 171018.245005086
Cbr48 netL48 0 -8.790590249832624e-21

* Branch 49
Rabr49 node_1 netRa49 48750.62595936208
Lbr49 netRa49 netL49 1.1413096323874179e-11
Rbbr49 netL49 0 -57514.53614566278
Cbr49 netL49 0 4.0715442292177974e-21

* Branch 50
Rabr50 node_1 netRa50 93062.51477168249
Lbr50 netRa50 netL50 1.0924519922408991e-10
Rbbr50 netL50 0 -399347.7897297749
Cbr50 netL50 0 2.9426172797303265e-21

* Branch 51
Rabr51 node_1 netRa51 558656.2329197116
Lbr51 netRa51 netL51 2.944499362367485e-10
Rbbr51 netL51 0 -783386.7269039764
Cbr51 netL51 0 6.731061210721674e-22

* Branch 52
Rabr52 node_1 netRa52 3853028.3422382385
Lbr52 netRa52 netL52 1.0481586117214655e-09
Rbbr52 netL52 0 -4162215.9711390412
Cbr52 netL52 0 6.537152731404687e-23

* Branch 53
Rabr53 node_1 netRa53 1976027.3418171594
Lbr53 netRa53 netL53 -3.236387124013632e-10
Rbbr53 netL53 0 -2090953.8992189667
Cbr53 netL53 0 -7.831997889034412e-23

* Branch 54
Rabr54 node_1 netRa54 113902.08769402986
Lbr54 netRa54 netL54 1.6398102307702575e-10
Rbbr54 netL54 0 -613700.1352836814
Cbr54 netL54 0 2.3478823412673165e-21

* Branch 55
Rabr55 node_1 netRa55 -316514.0055292932
Lbr55 netRa55 netL55 1.6488135770643859e-09
Rbbr55 netL55 0 17555917.32238756
Cbr55 netL55 0 2.9607142086016014e-22

* Branch 56
Rabr56 node_1 netRa56 -701123.0411552469
Lbr56 netRa56 netL56 -4.0747277690676396e-10
Rbbr56 netL56 0 1033527.2050915719
Cbr56 netL56 0 -5.624488641081247e-22

* Branch 57
Rabr57 node_1 netRa57 360493.23103499773
Lbr57 netRa57 netL57 8.925991561981686e-10
Rbbr57 netL57 0 -4055831.751976402
Cbr57 netL57 0 6.108624092678036e-22

* Branch 58
Rabr58 node_1 netRa58 -58584.44877876263
Lbr58 netRa58 netL58 -2.6677571034901945e-10
Rbbr58 netL58 0 1564914.0208758612
Cbr58 netL58 0 -2.9124420352914626e-21

* Branch 59
Rabr59 node_1 netRa59 -496735.40908145526
Lbr59 netRa59 netL59 7.844384284362218e-10
Rbbr59 netL59 0 2080988.8130846617
Cbr59 netL59 0 7.586621079117011e-22

* Branch 60
Rabr60 node_1 netRa60 361635.8353052218
Lbr60 netRa60 netL60 -1.4887368978766695e-10
Rbbr60 netL60 0 -442629.19215849537
Cbr60 netL60 0 -9.299905432592036e-22

* Branch 61
Rabr61 node_1 netRa61 343823.3449086273
Lbr61 netRa61 netL61 -7.039892242115344e-10
Rbbr61 netL61 0 -2554891.765740957
Cbr61 netL61 0 -8.012264657305349e-22

* Branch 62
Rabr62 node_1 netRa62 -11057290.070769517
Lbr62 netRa62 netL62 9.765373236471247e-09
Rbbr62 netL62 0 25868143.228492822
Cbr62 netL62 0 3.413757318320515e-23

* Branch 63
Rabr63 node_1 netRa63 10991239.725707365
Lbr63 netRa63 netL63 -1.4867865827050134e-09
Rbbr63 netL63 0 -11122613.977216255
Cbr63 netL63 0 -1.2161639442130704e-23

* Branch 64
Rabr64 node_1 netRa64 -65529.56340756273
Lbr64 netRa64 netL64 3.7462937466409233e-10
Rbbr64 netL64 0 911047.2119898791
Cbr64 netL64 0 6.274910681728908e-21

* Branch 65
Rabr65 node_1 netRa65 6530302.988616686
Lbr65 netRa65 netL65 -1.2570728955051016e-09
Rbbr65 netL65 0 -6757828.609118191
Cbr65 netL65 0 -2.848521121818366e-23

* Branch 66
Rabr66 node_1 netRa66 6176467.375682878
Lbr66 netRa66 netL66 -1.9628484605615066e-09
Rbbr66 netL66 0 -7337608.884628612
Cbr66 netL66 0 -4.3310304274708837e-23

* Branch 67
Rabr67 node_1 netRa67 2050980.9376406032
Lbr67 netRa67 netL67 -6.368229491998284e-10
Rbbr67 netL67 0 -2258082.9464497473
Cbr67 netL67 0 -1.3750277031624237e-22

* Branch 68
Rabr68 node_1 netRa68 363724.49102872994
Lbr68 netRa68 netL68 -3.610357717708614e-10
Rbbr68 netL68 0 -713216.8850232706
Cbr68 netL68 0 -1.391651306910962e-21

* Branch 69
Rabr69 node_1 netRa69 9352800.98316589
Lbr69 netRa69 netL69 1.8975243349146844e-09
Rbbr69 netL69 0 -9741976.550359152
Cbr69 netL69 0 2.0825917752976516e-23

* Branch 70
Rabr70 node_1 netRa70 1307154.0933939072
Lbr70 netRa70 netL70 -1.4799219813545932e-09
Rbbr70 netL70 0 -2352623.2662301334
Cbr70 netL70 0 -4.811962168775766e-22

* Branch 71
Rabr71 node_1 netRa71 2433487.363308051
Lbr71 netRa71 netL71 -6.972198753491343e-10
Rbbr71 netL71 0 -2795664.8863946423
Cbr71 netL71 0 -1.0248153957845658e-22

* Branch 72
Rabr72 node_1 netRa72 1990296.8812342188
Lbr72 netRa72 netL72 -1.0954894510150051e-09
Rbbr72 netL72 0 -2333179.140358726
Cbr72 netL72 0 -2.3589626448953846e-22

* Branch 73
Rabr73 node_1 netRa73 231189.26522749427
Lbr73 netRa73 netL73 -2.505784071302378e-10
Rbbr73 netL73 0 -378433.8817590787
Cbr73 netL73 0 -2.8638020292396887e-21

* Branch 74
Rabr74 node_1 netRa74 437952.4722351675
Lbr74 netRa74 netL74 -5.06974311765743e-10
Rbbr74 netL74 0 -787734.1764999484
Cbr74 netL74 0 -1.4693619799649309e-21

* Branch 75
Rabr75 node_1 netRa75 360677.6041120563
Lbr75 netRa75 netL75 -4.3360275072589956e-10
Rbbr75 netL75 0 -1207492.5427142966
Cbr75 netL75 0 -9.954582790889901e-22

* Branch 76
Rabr76 node_1 netRa76 528198.3875049466
Lbr76 netRa76 netL76 -5.37779407808674e-10
Rbbr76 netL76 0 -1494467.5629214344
Cbr76 netL76 0 -6.8118441392465635e-22

* Branch 77
Rabr77 node_1 netRa77 -2148852.708585978
Lbr77 netRa77 netL77 -1.0254814249709222e-09
Rbbr77 netL77 0 2735726.9588983473
Cbr77 netL77 0 -1.7445447198180675e-22

* Branch 78
Rabr78 node_1 netRa78 20580.208029808186
Lbr78 netRa78 netL78 -4.136689238031638e-10
Rbbr78 netL78 0 -3675059.6408230644
Cbr78 netL78 0 -5.446883406705408e-21

* Branch 79
Rabr79 node_1 netRa79 87232.81286877343
Lbr79 netRa79 netL79 6.109863391196991e-11
Rbbr79 netL79 0 -196672.49034649978
Cbr79 netL79 0 3.561860113943774e-21

* Branch 80
Rabr80 node_1 netRa80 5569929.865362174
Lbr80 netRa80 netL80 -7.14905418813785e-10
Rbbr80 netL80 0 -5778622.199106361
Cbr80 netL80 0 -2.2210644422556205e-23

* Branch 81
Rabr81 node_1 netRa81 77472.31227197054
Lbr81 netRa81 netL81 -2.7015565184296816e-10
Rbbr81 netL81 0 -1480376.1822768773
Cbr81 netL81 0 -2.3535590632019442e-21

* Branch 82
Rabr82 node_1 netRa82 76850.53043462327
Lbr82 netRa82 netL82 7.201880761596793e-11
Rbbr82 netL82 0 -168922.4951399578
Cbr82 netL82 0 5.549067581884204e-21

* Branch 83
Rabr83 node_1 netRa83 2132724.085353821
Lbr83 netRa83 netL83 4.5566115164543105e-10
Rbbr83 netL83 0 -2348936.362138941
Cbr83 netL83 0 9.096260874504686e-23

* Branch 84
Rabr84 node_1 netRa84 -1765692.4239919463
Lbr84 netRa84 netL84 -5.582029359366656e-10
Rbbr84 netL84 0 1970411.7189095756
Cbr84 netL84 0 -1.604579040695112e-22

* Branch 85
Rabr85 node_1 netRa85 126193.06861499159
Lbr85 netRa85 netL85 -1.399607518700548e-10
Rbbr85 netL85 0 -446312.07598437543
Cbr85 netL85 0 -2.4841570251865657e-21

* Branch 86
Rabr86 node_1 netRa86 82248.4235191142
Lbr86 netRa86 netL86 -8.540437718176072e-11
Rbbr86 netL86 0 -119441.26322267062
Cbr86 netL86 0 -8.690377949611375e-21

* Branch 87
Rabr87 node_1 netRa87 15665.108947236446
Lbr87 netRa87 netL87 3.51239932485683e-11
Rbbr87 netL87 0 -199500.29042559423
Cbr87 netL87 0 1.1248163660177521e-20

* Branch 88
Rabr88 node_1 netRa88 -4611.894095826369
Lbr88 netRa88 netL88 -1.1589162304938637e-10
Rbbr88 netL88 0 5779040.7585602235
Cbr88 netL88 0 -4.397038858159685e-21

* Branch 89
Rabr89 node_1 netRa89 32663.86335298063
Lbr89 netRa89 netL89 -1.3059098232367267e-10
Rbbr89 netL89 0 -419732.9558306711
Cbr89 netL89 0 -9.506896692647016e-21

* Branch 90
Rabr90 node_1 netRa90 123211.4810060218
Lbr90 netRa90 netL90 -2.8393890368945033e-10
Rbbr90 netL90 0 -629066.4111830115
Cbr90 netL90 0 -3.6587475321580306e-21

* Branch 91
Rabr91 node_1 netRa91 466141.9714499129
Lbr91 netRa91 netL91 -2.365931554697915e-10
Rbbr91 netL91 0 -551709.8447550775
Cbr91 netL91 0 -9.196735741641014e-22

* Branch 92
Rabr92 node_1 netRa92 87656.99362654924
Lbr92 netRa92 netL92 5.677060516091707e-11
Rbbr92 netL92 0 -194755.57384224495
Cbr92 netL92 0 3.3269381743173596e-21

* Branch 93
Rabr93 node_1 netRa93 95441.96935099683
Lbr93 netRa93 netL93 -9.725701965999768e-11
Rbbr93 netL93 0 -175282.57045609155
Cbr93 netL93 0 -5.809106250952137e-21

* Branch 94
Rabr94 node_1 netRa94 493984.5313804213
Lbr94 netRa94 netL94 8.668192016968509e-11
Rbbr94 netL94 0 -534629.4577800112
Cbr94 netL94 0 3.282664370725654e-22

* Branch 95
Rabr95 node_1 netRa95 -2591.9353300831285
Lbr95 netRa95 netL95 3.6229155156190678e-12
Rbbr95 netL95 0 18938.14673751032
Cbr95 netL95 0 7.368400364300867e-20

* Branch 96
Rabr96 node_1 netRa96 42218.09528572963
Lbr96 netRa96 netL96 2.905099666058375e-11
Rbbr96 netL96 0 -105464.2714198148
Cbr96 netL96 0 6.5302206088712314e-21

* Branch 97
Rabr97 node_1 netRa97 143680.6173203484
Lbr97 netRa97 netL97 3.873509240613896e-11
Rbbr97 netL97 0 -172222.04174404513
Cbr97 netL97 0 1.5659281706221555e-21

* Branch 98
Rabr98 node_1 netRa98 281565.17268607725
Lbr98 netRa98 netL98 -3.9054698433440936e-11
Rbbr98 netL98 0 -298357.4685079822
Cbr98 netL98 0 -4.647841464741996e-22

* Branch 99
Rabr99 node_1 netRa99 5824.106788088408
Lbr99 netRa99 netL99 -2.862532129830074e-12
Rbbr99 netL99 0 -10523.565209165967
Cbr99 netL99 0 -4.582883626100228e-20

.ends


* Y'12
.subckt yp12 node_1 node_2
* Branch 0
Rabr0 node_1 netRa0 -93.8986377214537
Lbr0 netRa0 netL0 1.306430107095016e-13
Rbbr0 netL0 node_2 377.0728025344691
Cbr0 netL0 node_2 3.153268525187051e-18

* Branch 1
Rabr1 node_1 netRa1 -40.10823038963884
Lbr1 netRa1 netL1 5.814250964792625e-14
Rbbr1 netL1 node_2 165.61115196748767
Cbr1 netL1 node_2 7.467001841788674e-18

* Branch 2
Rabr2 node_1 netRa2 -310.2950835823065
Lbr2 netRa2 netL2 1.4110856232680926e-13
Rbbr2 netL2 node_2 419.5065003231486
Cbr2 netL2 node_2 1.0370985642563338e-18

* Branch 3
Rabr3 node_1 netRa3 -487.6085384281788
Lbr3 netRa3 netL3 2.539536880613388e-13
Rbbr3 netL3 node_2 716.224866889084
Cbr3 netL3 node_2 6.927127870229529e-19

* Branch 4
Rabr4 node_1 netRa4 -2698.3712181840688
Lbr4 netRa4 netL4 4.089513821268382e-13
Rbbr4 netL4 node_2 2807.567133999856
Cbr4 netL4 node_2 5.3273593747816844e-20

* Branch 5
Rabr5 node_1 netRa5 153.49227831009682
Lbr5 netRa5 netL5 2.4460942973490186e-13
Rbbr5 netL5 node_2 -967.6391747458163
Cbr5 netL5 node_2 1.854796962181044e-18

* Branch 6
Rabr6 node_1 netRa6 66.07548835704554
Lbr6 netRa6 netL6 -3.56544792536057e-14
Rbbr6 netL6 node_2 -95.68804388247833
Cbr6 netL6 node_2 -5.449557384841234e-18

* Branch 7
Rabr7 node_1 netRa7 -26.543093408027815
Lbr7 netRa7 netL7 -7.655947193544539e-14
Rbbr7 netL7 node_2 486.68062255976264
Cbr7 netL7 node_2 -6.8359211183714775e-18

* Branch 8
Rabr8 node_1 netRa8 -5.587145496253745
Lbr8 netRa8 netL8 1.3563699853795534e-13
Rbbr8 netL8 node_2 2563.831585211404
Cbr8 netL8 node_2 4.751000849043171e-18

* Branch 9
Rabr9 node_1 netRa9 -112.25136786761517
Lbr9 netRa9 netL9 1.0827342955092167e-13
Rbbr9 netL9 node_2 268.6315660159456
Cbr9 netL9 node_2 3.4694306485485816e-18

* Branch 10
Rabr10 node_1 netRa10 -1202429.2891390962
Lbr10 netRa10 netL10 -1.1138649829740693e-11
Rbbr10 netL10 node_2 1202591.247015562
Cbr10 netL10 node_2 -7.705467879887805e-24

* Branch 11
Rabr11 node_1 netRa11 200.3258897914002
Lbr11 netRa11 netL11 7.570330209330387e-14
Rbbr11 netL11 node_2 -252.02064351305373
Cbr11 netL11 node_2 1.5196802646868807e-18

* Branch 12
Rabr12 node_1 netRa12 241.14733655182187
Lbr12 netRa12 netL12 -7.233230496932981e-14
Rbbr12 netL12 node_2 -280.4472289749641
Cbr12 netL12 node_2 -1.0586749421227908e-18

* Branch 13
Rabr13 node_1 netRa13 31998.956031408175
Lbr13 netRa13 netL13 -1.7153102195299182e-12
Rbbr13 netL13 node_2 -32156.25621803387
Cbr13 netL13 node_2 -1.663986989579704e-21

* Branch 14
Rabr14 node_1 netRa14 -70.29240821966471
Lbr14 netRa14 netL14 4.166317096708036e-14
Rbbr14 netL14 node_2 107.89985332041266
Cbr14 netL14 node_2 5.403728658187795e-18

* Branch 15
Rabr15 node_1 netRa15 140.38805395168555
Lbr15 netRa15 netL15 5.96352339231911e-14
Rbbr15 netL15 node_2 -180.67401240971233
Cbr15 netL15 node_2 2.3792793300086244e-18

* Branch 16
Rabr16 node_1 netRa16 -1885.5111515771498
Lbr16 netRa16 netL16 -5.809017049447567e-13
Rbbr16 netL16 node_2 2140.8356047984253
Cbr16 netL16 node_2 -1.451205444245278e-19

* Branch 17
Rabr17 node_1 netRa17 -6522.679533953477
Lbr17 netRa17 netL17 1.1709850663381918e-12
Rbbr17 netL17 node_2 6805.478747504596
Cbr17 netL17 node_2 2.6271712258744623e-20

* Branch 18
Rabr18 node_1 netRa18 -2221.887318626927
Lbr18 netRa18 netL18 -5.330899044149146e-13
Rbbr18 netL18 node_2 2410.505251547791
Cbr18 netL18 node_2 -1.0005433612488984e-19

* Branch 19
Rabr19 node_1 netRa19 -248.25095073721775
Lbr19 netRa19 netL19 2.260031792032255e-13
Rbbr19 netL19 node_2 878.2209613341126
Cbr19 netL19 node_2 1.0169044690881346e-18

* Branch 20
Rabr20 node_1 netRa20 -14217.947480682562
Lbr20 netRa20 netL20 1.6948560549261357e-12
Rbbr20 netL20 node_2 14833.055307445353
Cbr20 netL20 node_2 8.016297745376568e-21

* Branch 21
Rabr21 node_1 netRa21 -120073.79437596863
Lbr21 netRa21 netL21 1.2006300316272306e-11
Rbbr21 netL21 node_2 120635.72726181553
Cbr21 netL21 node_2 8.2718544920995e-22

* Branch 22
Rabr22 node_1 netRa22 -5588.050399164593
Lbr22 netRa22 netL22 1.4964274189325056e-12
Rbbr22 netL22 node_2 6871.179515697257
Cbr22 netL22 node_2 3.876924564518097e-20

* Branch 23
Rabr23 node_1 netRa23 -9450.770699658538
Lbr23 netRa23 netL23 -1.5379601987956191e-12
Rbbr23 netL23 node_2 10199.219781306578
Cbr23 netL23 node_2 -1.6005227189406777e-20

* Branch 24
Rabr24 node_1 netRa24 -218.60160610707592
Lbr24 netRa24 netL24 -1.29705055030079e-13
Rbbr24 netL24 node_2 336.5011268301105
Cbr24 netL24 node_2 -1.782679380101178e-18

* Branch 25
Rabr25 node_1 netRa25 8660.133747392798
Lbr25 netRa25 netL25 1.3448310289743306e-12
Rbbr25 netL25 node_2 -9360.25249452092
Cbr25 netL25 node_2 1.663762863466418e-20

* Branch 26
Rabr26 node_1 netRa26 33.34790901601987
Lbr26 netRa26 netL26 -5.97904098418687e-14
Rbbr26 netL26 node_2 -228.1197141117087
Cbr26 netL26 node_2 -7.613411057269939e-18

* Branch 27
Rabr27 node_1 netRa27 -2689.512228739211
Lbr27 netRa27 netL27 4.3878384834714316e-13
Rbbr27 netL27 node_2 2853.6011830639936
Cbr27 netL27 node_2 5.701321487250022e-20

* Branch 28
Rabr28 node_1 netRa28 604.3752742743923
Lbr28 netRa28 netL28 4.847558264109833e-13
Rbbr28 netL28 node_2 -1898.556077088233
Cbr28 netL28 node_2 4.278633301254332e-19

* Branch 29
Rabr29 node_1 netRa29 -489.6160184034313
Lbr29 netRa29 netL29 -4.24725750758165e-13
Rbbr29 netL29 node_2 804.2131046953035
Cbr29 netL29 node_2 -1.0918667088756362e-18

* Branch 30
Rabr30 node_1 netRa30 22870.504813394742
Lbr30 netRa30 netL30 -3.445187550709633e-12
Rbbr30 netL30 node_2 -24393.904427267826
Cbr30 netL30 node_2 -6.162755865593605e-21

* Branch 31
Rabr31 node_1 netRa31 -72190.89522175697
Lbr31 netRa31 netL31 3.675754437106337e-12
Rbbr31 netL31 node_2 72435.30115828967
Cbr31 netL31 node_2 7.024721479994876e-22

* Branch 32
Rabr32 node_1 netRa32 573.980259988249
Lbr32 netRa32 netL32 5.046469255732894e-13
Rbbr32 netL32 node_2 -1694.0561733846296
Cbr32 netL32 node_2 5.248559227299432e-19

* Branch 33
Rabr33 node_1 netRa33 -443.9729335267535
Lbr33 netRa33 netL33 -4.218361564088024e-13
Rbbr33 netL33 node_2 1627.2684518952826
Cbr33 netL33 node_2 -5.907862619341236e-19

* Branch 34
Rabr34 node_1 netRa34 9884.794544516353
Lbr34 netRa34 netL34 2.108974066820669e-12
Rbbr34 netL34 node_2 -11429.976296198589
Cbr34 netL34 node_2 1.8715330117372516e-20

* Branch 35
Rabr35 node_1 netRa35 -697.7788681839558
Lbr35 netRa35 netL35 1.9555923129356985e-13
Rbbr35 netL35 node_2 820.5356434472561
Cbr35 netL35 node_2 3.40390587509351e-19

* Branch 36
Rabr36 node_1 netRa36 -4533.145704781882
Lbr36 netRa36 netL36 8.126453963819391e-13
Rbbr36 netL36 node_2 4912.601735699819
Cbr36 netL36 node_2 3.641197557478616e-20

* Branch 37
Rabr37 node_1 netRa37 15.291892756564325
Lbr37 netRa37 netL37 -6.226373022777897e-14
Rbbr37 netL37 node_2 -316.15579875454813
Cbr37 netL37 node_2 -1.2332383292991816e-17

* Branch 38
Rabr38 node_1 netRa38 15841.346801408901
Lbr38 netRa38 netL38 2.2763120732135573e-12
Rbbr38 netL38 node_2 -16895.601002879383
Cbr38 netL38 node_2 8.516664871643869e-21

* Branch 39
Rabr39 node_1 netRa39 -163.6469849347797
Lbr39 netRa39 netL39 -2.2766158350958366e-13
Rbbr39 netL39 node_2 458.4878119108506
Cbr39 netL39 node_2 -3.0744049341959714e-18

* Branch 40
Rabr40 node_1 netRa40 16.184677267314818
Lbr40 netRa40 netL40 -1.2017073050149982e-13
Rbbr40 netL40 node_2 -988.1477058755431
Cbr40 netL40 node_2 -7.05185583278786e-18

* Branch 41
Rabr41 node_1 netRa41 1030.2715458297764
Lbr41 netRa41 netL41 4.894836097071469e-13
Rbbr41 netL41 node_2 -1597.3965457047066
Cbr41 netL41 node_2 2.9867475967543567e-19

* Branch 42
Rabr42 node_1 netRa42 3119.0844697803136
Lbr42 netRa42 netL42 1.0873296984351756e-12
Rbbr42 netL42 node_2 -4319.72331894191
Cbr42 netL42 node_2 8.093784487258084e-20

* Branch 43
Rabr43 node_1 netRa43 -644.4289755963391
Lbr43 netRa43 netL43 -5.387198767787022e-13
Rbbr43 netL43 node_2 985.8190933919881
Cbr43 netL43 node_2 -8.539478226986535e-19

* Branch 44
Rabr44 node_1 netRa44 92009.1377968801
Lbr44 netRa44 netL44 6.3728647538202116e-12
Rbbr44 netL44 node_2 -93136.22422238666
Cbr44 netL44 node_2 7.440721112044843e-22

* Branch 45
Rabr45 node_1 netRa45 -69.51679249921384
Lbr45 netRa45 netL45 -1.5964974818223396e-13
Rbbr45 netL45 node_2 442.2481267311618
Cbr45 netL45 node_2 -5.274740039526268e-18

* Branch 46
Rabr46 node_1 netRa46 718.5639586308291
Lbr46 netRa46 netL46 5.051334724988281e-13
Rbbr46 netL46 node_2 -1668.396390500857
Cbr46 netL46 node_2 4.231998896471914e-19

* Branch 47
Rabr47 node_1 netRa47 12842.896947687694
Lbr47 netRa47 netL47 3.011951559494564e-12
Rbbr47 netL47 node_2 -15312.43603743136
Cbr47 netL47 node_2 1.5337036991010094e-20

* Branch 48
Rabr48 node_1 netRa48 13.055617484470222
Lbr48 netRa48 netL48 -1.8269001703605864e-13
Rbbr48 netL48 node_2 -4536.418646138366
Cbr48 netL48 node_2 -2.850683097909374e-18

* Branch 49
Rabr49 node_1 netRa49 -639.1116797133337
Lbr49 netRa49 netL49 -2.980016653189777e-13
Rbbr49 netL49 node_2 938.6399386822728
Cbr49 netL49 node_2 -4.980516207894649e-19

* Branch 50
Rabr50 node_1 netRa50 -1302.7899845754823
Lbr50 netRa50 netL50 2.920088230884707e-13
Rbbr50 netL50 node_2 1455.467624332698
Cbr50 netL50 node_2 1.5380994573821576e-19

* Branch 51
Rabr51 node_1 netRa51 -6699.32344133412
Lbr51 netRa51 netL51 -2.025370786088076e-12
Rbbr51 netL51 node_2 7115.82445108944
Cbr51 netL51 node_2 -4.255279162845768e-20

* Branch 52
Rabr52 node_1 netRa52 -328.4750283775336
Lbr52 netRa52 netL52 -4.685156468242834e-13
Rbbr52 netL52 node_2 2114.772674797393
Cbr52 netL52 node_2 -6.793997232329062e-19

* Branch 53
Rabr53 node_1 netRa53 -34472216.735019565
Lbr53 netRa53 netL53 1.806496385296116e-10
Rbbr53 netL53 node_2 34472729.99197607
Cbr53 netL53 node_2 1.5201312498874143e-25

* Branch 54
Rabr54 node_1 netRa54 -593.6014551012836
Lbr54 netRa54 netL54 -2.2676272017643363e-13
Rbbr54 netL54 node_2 774.9656249759894
Cbr54 netL54 node_2 -4.937683035448074e-19

* Branch 55
Rabr55 node_1 netRa55 4463.916123402828
Lbr55 netRa55 netL55 -1.5109318617148002e-12
Rbbr55 netL55 node_2 -5882.62730046013
Cbr55 netL55 node_2 -5.747740777952875e-20

* Branch 56
Rabr56 node_1 netRa56 2513.4686038377613
Lbr56 netRa56 netL56 5.66578942536464e-13
Rbbr56 netL56 node_2 -2816.83612896378
Cbr56 netL56 node_2 8.007936786196872e-20

* Branch 57
Rabr57 node_1 netRa57 -133.55230301435714
Lbr57 netRa57 netL57 3.2274116267318575e-13
Rbbr57 netL57 node_2 1033.260413627482
Cbr57 netL57 node_2 2.322271191159401e-18

* Branch 58
Rabr58 node_1 netRa58 1624.2872148278334
Lbr58 netRa58 netL58 -1.0266728062782458e-12
Rbbr58 netL58 node_2 -3461.4487909346703
Cbr58 netL58 node_2 -1.8226606401345246e-19

* Branch 59
Rabr59 node_1 netRa59 -704.5812378046343
Lbr59 netRa59 netL59 -2.94701659887218e-13
Rbbr59 netL59 node_2 976.8513152456222
Cbr59 netL59 node_2 -4.286765378276524e-19

* Branch 60
Rabr60 node_1 netRa60 356721.22704296495
Lbr60 netRa60 netL60 -2.41425290613936e-11
Rbbr60 netL60 node_2 -358552.07376480015
Cbr60 netL60 node_2 -1.8872613686423062e-22

* Branch 61
Rabr61 node_1 netRa61 404.25035487689087
Lbr61 netRa61 netL61 -3.7291512810675664e-13
Rbbr61 netL61 node_2 -1183.1185973067345
Cbr61 netL61 node_2 -7.780612084634129e-19

* Branch 62
Rabr62 node_1 netRa62 1499.418837670276
Lbr62 netRa62 netL62 -8.709314719167949e-13
Rbbr62 netL62 node_2 -2816.3863227935476
Cbr62 netL62 node_2 -2.0597431665157672e-19

* Branch 63
Rabr63 node_1 netRa63 6423.97529823755
Lbr63 netRa63 netL63 5.579014098823113e-12
Rbbr63 netL63 node_2 -10181.310232170163
Cbr63 netL63 node_2 8.545130601746598e-20

* Branch 64
Rabr64 node_1 netRa64 4795.170206233212
Lbr64 netRa64 netL64 -1.7693889351886102e-12
Rbbr64 netL64 node_2 -6570.2818219621495
Cbr64 netL64 node_2 -5.611909407657878e-20

* Branch 65
Rabr65 node_1 netRa65 6471.506712252993
Lbr65 netRa65 netL65 -5.33742815674815e-12
Rbbr65 netL65 node_2 -9213.482661392709
Cbr65 netL65 node_2 -8.937510004957676e-20

* Branch 66
Rabr66 node_1 netRa66 901.2282377896128
Lbr66 netRa66 netL66 1.3413439189971437e-12
Rbbr66 netL66 node_2 -8035.136940131702
Cbr66 netL66 node_2 1.857531972471539e-19

* Branch 67
Rabr67 node_1 netRa67 46132.69658952534
Lbr67 netRa67 netL67 1.2743358427465036e-11
Rbbr67 netL67 node_2 -48972.27706273204
Cbr67 netL67 node_2 5.642759708740402e-21

* Branch 68
Rabr68 node_1 netRa68 -50.11031418303911
Lbr68 netRa68 netL68 -1.7010480739731476e-13
Rbbr68 netL68 node_2 1396.5702907557152
Cbr68 netL68 node_2 -2.4420749036581735e-18

* Branch 69
Rabr69 node_1 netRa69 -2726.4613595164333
Lbr69 netRa69 netL69 5.320565657451467e-12
Rbbr69 netL69 node_2 13579.922174643134
Cbr69 netL69 node_2 1.4332480998051213e-19

* Branch 70
Rabr70 node_1 netRa70 3814.4304646518012
Lbr70 netRa70 netL70 6.408707235756872e-12
Rbbr70 netL70 node_2 -15519.523935966272
Cbr70 netL70 node_2 1.0849055990581173e-19

* Branch 71
Rabr71 node_1 netRa71 392.48619301224727
Lbr71 netRa71 netL71 5.134672024053171e-13
Rbbr71 netL71 node_2 -1224.9737220575964
Cbr71 netL71 node_2 1.069525206700561e-18

* Branch 72
Rabr72 node_1 netRa72 48088.59253166986
Lbr72 netRa72 netL72 -1.664705003150549e-11
Rbbr72 netL72 node_2 -51516.069037102454
Cbr72 netL72 node_2 -6.717247915979904e-21

* Branch 73
Rabr73 node_1 netRa73 -3210.483078740621
Lbr73 netRa73 netL73 1.8673666782845836e-12
Rbbr73 netL73 node_2 4596.380590442511
Cbr73 netL73 node_2 1.2647629180032357e-19

* Branch 74
Rabr74 node_1 netRa74 9871.346873698036
Lbr74 netRa74 netL74 -5.344977761061234e-12
Rbbr74 netL74 node_2 -12295.040398193903
Cbr74 netL74 node_2 -4.4018870354792666e-20

* Branch 75
Rabr75 node_1 netRa75 -3938.406966348624
Lbr75 netRa75 netL75 -1.2487907262073394e-12
Rbbr75 netL75 node_2 4713.74019168377
Cbr75 netL75 node_2 -6.728519560700679e-20

* Branch 76
Rabr76 node_1 netRa76 -1470.467249819343
Lbr76 netRa76 netL76 2.398386675999007e-12
Rbbr76 netL76 node_2 5419.61915023118
Cbr76 netL76 node_2 3.0054825741228083e-19

* Branch 77
Rabr77 node_1 netRa77 1741.802155075948
Lbr77 netRa77 netL77 4.5915077785366535e-12
Rbbr77 netL77 node_2 -16287.164737895999
Cbr77 netL77 node_2 1.6214900347716302e-19

* Branch 78
Rabr78 node_1 netRa78 -5084.830336330507
Lbr78 netRa78 netL78 4.995243441278929e-12
Rbbr78 netL78 node_2 9700.018655797909
Cbr78 netL78 node_2 1.0122048761219218e-19

* Branch 79
Rabr79 node_1 netRa79 1601.755671884928
Lbr79 netRa79 netL79 3.9871812304618165e-12
Rbbr79 netL79 node_2 -11297.652826880167
Cbr79 netL79 node_2 2.2060491680906106e-19

* Branch 80
Rabr80 node_1 netRa80 -3210.4250885843758
Lbr80 netRa80 netL80 -1.6444280247537312e-12
Rbbr80 netL80 node_2 3704.5498681918216
Cbr80 netL80 node_2 -1.382889705173981e-19

* Branch 81
Rabr81 node_1 netRa81 9792.175804181998
Lbr81 netRa81 netL81 8.901424829566626e-12
Rbbr81 netL81 node_2 -17121.536942733368
Cbr81 netL81 node_2 5.310705629263256e-20

* Branch 82
Rabr82 node_1 netRa82 558.823138126166
Lbr82 netRa82 netL82 -7.443614928949544e-12
Rbbr82 netL82 node_2 -65004.477574692755
Cbr82 netL82 node_2 -2.041992279126383e-19

* Branch 83
Rabr83 node_1 netRa83 65205.9596273438
Lbr83 netRa83 netL83 -3.2554874371229427e-11
Rbbr83 netL83 node_2 -79365.84951822674
Cbr83 netL83 node_2 -6.289888412513695e-21

* Branch 84
Rabr84 node_1 netRa84 2480.5980291685814
Lbr84 netRa84 netL84 -9.844551526058841e-12
Rbbr84 netL84 node_2 -30258.141373092345
Cbr84 netL84 node_2 -1.3105051042325353e-19

* Branch 85
Rabr85 node_1 netRa85 -213.48082901875418
Lbr85 netRa85 netL85 -3.187117896690335e-12
Rbbr85 netL85 node_2 35580.33100826631
Cbr85 netL85 node_2 -4.2039992169089844e-19

* Branch 86
Rabr86 node_1 netRa86 899.6663494487696
Lbr86 netRa86 netL86 -2.062952916460744e-12
Rbbr86 netL86 node_2 -4120.512521240618
Cbr86 netL86 node_2 -5.56411148804452e-19

* Branch 87
Rabr87 node_1 netRa87 -1876.240761270377
Lbr87 netRa87 netL87 -8.162905177670624e-12
Rbbr87 netL87 node_2 16695.65472203734
Cbr87 netL87 node_2 -2.606322352406049e-19

* Branch 88
Rabr88 node_1 netRa88 -4428.939220275832
Lbr88 netRa88 netL88 -1.8317252821257862e-11
Rbbr88 netL88 node_2 43481.40527047479
Cbr88 netL88 node_2 -9.512879810041535e-20

* Branch 89
Rabr89 node_1 netRa89 577.7125527847238
Lbr89 netRa89 netL89 -5.625702646480074e-13
Rbbr89 netL89 node_2 -2164.255550675746
Cbr89 netL89 node_2 -4.499341588208415e-19

* Branch 90
Rabr90 node_1 netRa90 -1700.4767543336739
Lbr90 netRa90 netL90 -6.906604551704971e-12
Rbbr90 netL90 node_2 14063.20108485826
Cbr90 netL90 node_2 -2.8881172092182798e-19

* Branch 91
Rabr91 node_1 netRa91 -467.1438803539255
Lbr91 netRa91 netL91 -6.090844840478353e-12
Rbbr91 netL91 node_2 39363.061213456625
Cbr91 netL91 node_2 -3.3134918827512174e-19

* Branch 92
Rabr92 node_1 netRa92 -474.52335718445903
Lbr92 netRa92 netL92 -4.311397165299823e-12
Rbbr92 netL92 node_2 18691.85363264412
Cbr92 netL92 node_2 -4.863345171890973e-19

* Branch 93
Rabr93 node_1 netRa93 -319.0204766478155
Lbr93 netRa93 netL93 -7.816485532175029e-12
Rbbr93 netL93 node_2 109307.13451733811
Cbr93 netL93 node_2 -2.2455902121892414e-19

* Branch 94
Rabr94 node_1 netRa94 365.04132773251564
Lbr94 netRa94 netL94 -2.6436503674246627e-12
Rbbr94 netL94 node_2 -10705.207557189022
Cbr94 netL94 node_2 -6.751013813124622e-19

* Branch 95
Rabr95 node_1 netRa95 1962.0231521403625
Lbr95 netRa95 netL95 4.819763439335218e-12
Rbbr95 netL95 node_2 -6640.075929114415
Cbr95 netL95 node_2 3.702944499569561e-19

* Branch 96
Rabr96 node_1 netRa96 -804.2733425062139
Lbr96 netRa96 netL96 -7.270807745301785e-13
Rbbr96 netL96 node_2 2125.25235957884
Cbr96 netL96 node_2 -4.255826597733721e-19

* Branch 97
Rabr97 node_1 netRa97 -115.92094034131071
Lbr97 netRa97 netL97 -1.2709805957420538e-13
Rbbr97 netL97 node_2 403.1082663330855
Cbr97 netL97 node_2 -2.733974435203627e-18

* Branch 98
Rabr98 node_1 netRa98 642.5135406507079
Lbr98 netRa98 netL98 -2.1965759634088775e-13
Rbbr98 netL98 node_2 -757.2034031509742
Cbr98 netL98 node_2 -4.429798445382821e-19

* Branch 99
Rabr99 node_1 netRa99 -137.18843880028732
Lbr99 netRa99 netL99 9.83395680744528e-14
Rbbr99 netL99 node_2 253.12643511456662
Cbr99 netL99 node_2 2.6275639786255126e-18

.ends


* Y'13
.subckt yp13 node_1 node_3
* Branch 0
Rabr0 node_1 netRa0 -57154.1890557577
Lbr0 netRa0 netL0 1.2472396451378826e-11
Rbbr0 netL0 node_3 64566.91254290912
Cbr0 netL0 node_3 3.3535495658099484e-21

* Branch 1
Rabr1 node_1 netRa1 -113.38036925534239
Lbr1 netRa1 netL1 -3.841009380194765e-12
Rbbr1 netL1 node_3 5638687.437582718
Cbr1 netL1 node_3 -9.453181763316509e-20

* Branch 2
Rabr2 node_1 netRa2 -1534.998367959483
Lbr2 netRa2 netL2 1.6224034766102303e-12
Rbbr2 netL2 node_3 6839.512421510858
Cbr2 netL2 node_3 1.5053029708435381e-19

* Branch 3
Rabr3 node_1 netRa3 -431.4340658203595
Lbr3 netRa3 netL3 1.94045793895313e-12
Rbbr3 netL3 node_3 20399.241585188727
Cbr3 netL3 node_3 1.9843252632380752e-19

* Branch 4
Rabr4 node_1 netRa4 -98.40226857661067
Lbr4 netRa4 netL4 4.768387600833346e-12
Rbbr4 netL4 node_3 196774.19201739496
Cbr4 netL4 node_3 1.1553489572472038e-19

* Branch 5
Rabr5 node_1 netRa5 -270.2842190461722
Lbr5 netRa5 netL5 -2.331648646527936e-12
Rbbr5 netL5 node_3 74486.92749649943
Cbr5 netL5 node_3 -1.4320512293866477e-19

* Branch 6
Rabr6 node_1 netRa6 18853.934458931995
Lbr6 netRa6 netL6 -3.754081519116397e-12
Rbbr6 netL6 node_3 -20913.116173979066
Cbr6 netL6 node_3 -9.479957868194981e-21

* Branch 7
Rabr7 node_1 netRa7 1459.0695999167706
Lbr7 netRa7 netL7 3.3672636852837134e-12
Rbbr7 netL7 node_3 -18256.90415691392
Cbr7 netL7 node_3 1.3303640316940592e-19

* Branch 8
Rabr8 node_1 netRa8 -137908.98802196365
Lbr8 netRa8 netL8 -1.191411673305937e-11
Rbbr8 netL8 node_3 140872.71346514145
Cbr8 netL8 node_3 -6.143658521441191e-22

* Branch 9
Rabr9 node_1 netRa9 2078.282034339947
Lbr9 netRa9 netL9 3.091343392038065e-12
Rbbr9 netL9 node_3 -13062.094570398503
Cbr9 netL9 node_3 1.174542174792074e-19

* Branch 10
Rabr10 node_1 netRa10 47747.564159451875
Lbr10 netRa10 netL10 -2.8122717785206295e-11
Rbbr10 netL10 node_3 -78593.34113052428
Cbr10 netL10 node_3 -7.405768939516052e-21

* Branch 11
Rabr11 node_1 netRa11 -993.9011991230108
Lbr11 netRa11 netL11 9.366900188126346e-13
Rbbr11 netL11 node_3 3430.7921054547874
Cbr11 netL11 node_3 2.6958615864914447e-19

* Branch 12
Rabr12 node_1 netRa12 -40893.15015488229
Lbr12 netRa12 netL12 1.253769026283993e-11
Rbbr12 netL12 node_3 52600.55148801429
Cbr12 netL12 node_3 5.7937504408059614e-21

* Branch 13
Rabr13 node_1 netRa13 2820.591263335119
Lbr13 netRa13 netL13 5.052045516549742e-12
Rbbr13 netL13 node_3 -23609.633705901106
Cbr13 netL13 node_3 7.849083248661418e-20

* Branch 14
Rabr14 node_1 netRa14 8431.439949517064
Lbr14 netRa14 netL14 2.443035657061834e-12
Rbbr14 netL14 node_3 -10295.548830031761
Cbr14 netL14 node_3 2.8292520926068157e-20

* Branch 15
Rabr15 node_1 netRa15 677.2213278886663
Lbr15 netRa15 netL15 1.0520810458005293e-11
Rbbr15 netL15 node_3 -395524.00789192825
Cbr15 netL15 node_3 5.443498805079643e-20

* Branch 16
Rabr16 node_1 netRa16 -932.487594030062
Lbr16 netRa16 netL16 8.553320825491232e-13
Rbbr16 netL16 node_3 3024.9585854794595
Cbr16 netL16 node_3 2.984076704038728e-19

* Branch 17
Rabr17 node_1 netRa17 10402.594162695641
Lbr17 netRa17 netL17 1.8538585848338596e-11
Rbbr17 netL17 node_3 -59437.86103546724
Cbr17 netL17 node_3 3.094699104602784e-20

* Branch 18
Rabr18 node_1 netRa18 174.31241984934897
Lbr18 netRa18 netL18 3.699147010459283e-12
Rbbr18 netL18 node_3 -155239.7854958253
Cbr18 netL18 node_3 2.0997589140378782e-19

* Branch 19
Rabr19 node_1 netRa19 51.10575271209643
Lbr19 netRa19 netL19 3.541801462907943e-12
Rbbr19 netL19 node_3 3165172.869483644
Cbr19 netL19 node_3 1.6635507496863534e-19

* Branch 20
Rabr20 node_1 netRa20 6380.594899157172
Lbr20 netRa20 netL20 8.392298526913724e-12
Rbbr20 netL20 node_3 -23669.626926374833
Cbr20 netL20 node_3 5.672718883564557e-20

* Branch 21
Rabr21 node_1 netRa21 -93488.30323126198
Lbr21 netRa21 netL21 2.6440347624593076e-11
Rbbr21 netL21 node_3 103411.85825053167
Cbr21 netL21 node_3 2.7231709295344558e-21

* Branch 22
Rabr22 node_1 netRa22 -2737.6989172795397
Lbr22 netRa22 netL22 6.989334835976357e-12
Rbbr22 netL22 node_3 26799.459247658455
Cbr22 netL22 node_3 9.172980066362876e-20

* Branch 23
Rabr23 node_1 netRa23 -19932.200932674517
Lbr23 netRa23 netL23 7.48300359651591e-12
Rbbr23 netL23 node_3 25987.58813599175
Cbr23 netL23 node_3 1.4365422409209656e-20

* Branch 24
Rabr24 node_1 netRa24 -217.8283891964092
Lbr24 netRa24 netL24 2.2379602647661365e-12
Rbbr24 netL24 node_3 66006.58830826789
Cbr24 netL24 node_3 1.350040728635067e-19

* Branch 25
Rabr25 node_1 netRa25 3439.1809965117
Lbr25 netRa25 netL25 6.328925365015312e-12
Rbbr25 netL25 node_3 -22445.633042828154
Cbr25 netL25 node_3 8.419342167826328e-20

* Branch 26
Rabr26 node_1 netRa26 -339420.5793457955
Lbr26 netRa26 netL26 -3.935993515800199e-11
Rbbr26 netL26 node_3 354394.22137758636
Cbr26 netL26 node_3 -3.2774562464029464e-22

* Branch 27
Rabr27 node_1 netRa27 -4133840.8773080823
Lbr27 netRa27 netL27 1.33138144718377e-10
Rbbr27 netL27 node_3 4142904.20130614
Cbr27 netL27 node_3 7.770702510645649e-24

* Branch 28
Rabr28 node_1 netRa28 -755.7321913640676
Lbr28 netRa28 netL28 1.1952122126308708e-12
Rbbr28 netL28 node_3 5283.725802774675
Cbr28 netL28 node_3 2.9361774401396136e-19

* Branch 29
Rabr29 node_1 netRa29 2654.1746423180134
Lbr29 netRa29 netL29 6.077146884667428e-12
Rbbr29 netL29 node_3 -18938.528621364763
Cbr29 netL29 node_3 1.243596268322809e-19

* Branch 30
Rabr30 node_1 netRa30 -10941.633774583937
Lbr30 netRa30 netL30 9.683133226071112e-12
Rbbr30 netL30 node_3 22444.329594180304
Cbr30 netL30 node_3 3.9014827083936765e-20

* Branch 31
Rabr31 node_1 netRa31 5696.896551373293
Lbr31 netRa31 netL31 8.855302714632634e-12
Rbbr31 netL31 node_3 -20272.06359388997
Cbr31 netL31 node_3 7.806781243857952e-20

* Branch 32
Rabr32 node_1 netRa32 2221.684896958872
Lbr32 netRa32 netL32 6.05248350507858e-12
Rbbr32 netL32 node_3 -17057.45625567771
Cbr32 netL32 node_3 1.643851578197674e-19

* Branch 33
Rabr33 node_1 netRa33 6293.407657104197
Lbr33 netRa33 netL33 1.0928081776971197e-11
Rbbr33 netL33 node_3 -20680.155312641084
Cbr33 netL33 node_3 8.548294778328345e-20

* Branch 34
Rabr34 node_1 netRa34 24651.18935154252
Lbr34 netRa34 netL34 2.5525568264985124e-11
Rbbr34 netL34 node_3 -39674.72234862433
Cbr34 netL34 node_3 2.637347675132636e-20

* Branch 35
Rabr35 node_1 netRa35 -15352.87469552815
Lbr35 netRa35 netL35 2.143787641755334e-11
Rbbr35 netL35 node_3 42441.54782758737
Cbr35 netL35 node_3 3.245083155584292e-20

* Branch 36
Rabr36 node_1 netRa36 17357.488648144845
Lbr36 netRa36 netL36 8.258524264283194e-12
Rbbr36 netL36 node_3 -25106.44654916034
Cbr36 netL36 node_3 1.904035903168362e-20

* Branch 37
Rabr37 node_1 netRa37 -121851.17884178115
Lbr37 netRa37 netL37 -2.2656819936836875e-11
Rbbr37 netL37 node_3 135163.09419314348
Cbr37 netL37 node_3 -1.3777986731596749e-21

* Branch 38
Rabr38 node_1 netRa38 2240.7119443721226
Lbr38 netRa38 netL38 3.873522269475244e-12
Rbbr38 netL38 node_3 -25480.28552806596
Cbr38 netL38 node_3 6.881942192885419e-20

* Branch 39
Rabr39 node_1 netRa39 -12262.026380470577
Lbr39 netRa39 netL39 6.46886824718549e-12
Rbbr39 netL39 node_3 24030.380141927337
Cbr39 netL39 node_3 2.186374843300662e-20

* Branch 40
Rabr40 node_1 netRa40 4648.473780777855
Lbr40 netRa40 netL40 8.818051951607533e-12
Rbbr40 netL40 node_3 -18426.413821879807
Cbr40 netL40 node_3 1.0438907062040563e-19

* Branch 41
Rabr41 node_1 netRa41 13666.63874867532
Lbr41 netRa41 netL41 1.809670266379757e-11
Rbbr41 netL41 node_3 -28099.5427369208
Cbr41 netL41 node_3 4.7577845206237524e-20

* Branch 42
Rabr42 node_1 netRa42 651884.0457679849
Lbr42 netRa42 netL42 2.3261348691716842e-11
Rbbr42 netL42 node_3 -654326.5208598013
Cbr42 netL42 node_3 5.454651576382493e-23

* Branch 43
Rabr43 node_1 netRa43 8238.08389135336
Lbr43 netRa43 netL43 1.084958151848246e-11
Rbbr43 netL43 node_3 -22517.146590498633
Cbr43 netL43 node_3 5.895792259969635e-20

* Branch 44
Rabr44 node_1 netRa44 -168943.6258229139
Lbr44 netRa44 netL44 -5.3327085935808894e-11
Rbbr44 netL44 node_3 184794.6706802743
Cbr44 netL44 node_3 -1.7107308820174034e-21

* Branch 45
Rabr45 node_1 netRa45 3951.2546248787035
Lbr45 netRa45 netL45 -7.191631812252407e-12
Rbbr45 netL45 node_3 -9669.224142795563
Cbr45 netL45 node_3 -1.8675495233078824e-19

* Branch 46
Rabr46 node_1 netRa46 -7211.130543403791
Lbr46 netRa46 netL46 -1.7048689407179328e-11
Rbbr46 netL46 node_3 28322.908516685424
Cbr46 netL46 node_3 -8.41904162102835e-20

* Branch 47
Rabr47 node_1 netRa47 -664.8708179134245
Lbr47 netRa47 netL47 -2.4517839157803235e-11
Rbbr47 netL47 node_3 510468.9331102329
Cbr47 netL47 node_3 -8.301062868211898e-20

* Branch 48
Rabr48 node_1 netRa48 -6617.12998269671
Lbr48 netRa48 netL48 1.3188066456362543e-11
Rbbr48 netL48 node_3 50187.04176417169
Cbr48 netL48 node_3 3.944368038830964e-20

* Branch 49
Rabr49 node_1 netRa49 282.35091459481123
Lbr49 netRa49 netL49 1.1903496841929533e-11
Rbbr49 netL49 node_3 -703214.2407552375
Cbr49 netL49 node_3 6.996560446748029e-20

* Branch 50
Rabr50 node_1 netRa50 -16786.129694582873
Lbr50 netRa50 netL50 1.6005308669461e-11
Rbbr50 netL50 node_3 41461.50164615144
Cbr50 netL50 node_3 2.2923005489864484e-20

* Branch 51
Rabr51 node_1 netRa51 506.24056812872067
Lbr51 netRa51 netL51 -2.0261953758578652e-12
Rbbr51 netL51 node_3 -21996.078852145038
Cbr51 netL51 node_3 -1.796011714799556e-19

* Branch 52
Rabr52 node_1 netRa52 -10710.729188888185
Lbr52 netRa52 netL52 -6.658174157361591e-12
Rbbr52 netL52 node_3 19960.5204452657
Cbr52 netL52 node_3 -3.1204382117938695e-20

* Branch 53
Rabr53 node_1 netRa53 7813.253314557401
Lbr53 netRa53 netL53 1.3256433024125951e-11
Rbbr53 netL53 node_3 -22791.79723929345
Cbr53 netL53 node_3 7.477887770970011e-20

* Branch 54
Rabr54 node_1 netRa54 115126.49535583064
Lbr54 netRa54 netL54 -1.644102626920977e-11
Rbbr54 netL54 node_3 -121799.36658445098
Cbr54 netL54 node_3 -1.1721027510808356e-21

* Branch 55
Rabr55 node_1 netRa55 -2631.7300952905857
Lbr55 netRa55 netL55 1.0574213995833388e-11
Rbbr55 netL55 node_3 83260.71737424153
Cbr55 netL55 node_3 4.7892981505826355e-20

* Branch 56
Rabr56 node_1 netRa56 2748.596784896699
Lbr56 netRa56 netL56 1.820800168550743e-11
Rbbr56 netL56 node_3 -144304.64100036724
Cbr56 netL56 node_3 4.643719565668133e-20

* Branch 57
Rabr57 node_1 netRa57 -710.1267831839605
Lbr57 netRa57 netL57 1.2545016577631225e-11
Rbbr57 netL57 node_3 502392.63583740353
Cbr57 netL57 node_3 3.417765409128053e-20

* Branch 58
Rabr58 node_1 netRa58 -58527.60256204557
Lbr58 netRa58 netL58 2.2925489813470526e-11
Rbbr58 netL58 node_3 79910.04981379276
Cbr58 netL58 node_3 4.898748773495658e-21

* Branch 59
Rabr59 node_1 netRa59 -229225.6602586662
Lbr59 netRa59 netL59 5.424781236713192e-11
Rbbr59 netL59 node_3 270601.59708684863
Cbr59 netL59 node_3 8.742282544513775e-22

* Branch 60
Rabr60 node_1 netRa60 -19402.013077740066
Lbr60 netRa60 netL60 1.696175923020183e-11
Rbbr60 netL60 node_3 40890.0391773426
Cbr60 netL60 node_3 2.1352224822974984e-20

* Branch 61
Rabr61 node_1 netRa61 -1328.846285852195
Lbr61 netRa61 netL61 8.677530067205724e-12
Rbbr61 netL61 node_3 116975.0318419298
Cbr61 netL61 node_3 5.533611152673064e-20

* Branch 62
Rabr62 node_1 netRa62 -4259617.171904152
Lbr62 netRa62 netL62 2.1724617332510083e-10
Rbbr62 netL62 node_3 4279176.816555884
Cbr62 netL62 node_3 1.1917948032923467e-23

* Branch 63
Rabr63 node_1 netRa63 -1277.0658455703956
Lbr63 netRa63 netL63 1.4244031775299836e-11
Rbbr63 netL63 node_3 317997.70095993945
Cbr63 netL63 node_3 3.479399125378461e-20

* Branch 64
Rabr64 node_1 netRa64 -375810.93368732324
Lbr64 netRa64 netL64 1.0567586454963429e-10
Rbbr64 netL64 node_3 420093.8536113393
Cbr64 netL64 node_3 6.692334386434719e-22

* Branch 65
Rabr65 node_1 netRa65 11889.884851664912
Lbr65 netRa65 netL65 3.290179209460124e-11
Rbbr65 netL65 node_3 -74035.22611695672
Cbr65 netL65 node_3 3.743641322722151e-20

* Branch 66
Rabr66 node_1 netRa66 6412.1327759818
Lbr66 netRa66 netL66 3.124180614901768e-11
Rbbr66 netL66 node_3 -160527.32095362773
Cbr66 netL66 node_3 3.041519121690168e-20

* Branch 67
Rabr67 node_1 netRa67 12873.351269663268
Lbr67 netRa67 netL67 3.440096794218161e-11
Rbbr67 netL67 node_3 -78350.3682660702
Cbr67 netL67 node_3 3.4143356005611165e-20

* Branch 68
Rabr68 node_1 netRa68 -71573.14448668616
Lbr68 netRa68 netL68 4.607750528335734e-11
Rbbr68 netL68 node_3 125334.0672190955
Cbr68 netL68 node_3 5.1352950586257555e-21

* Branch 69
Rabr69 node_1 netRa69 15414.584429316868
Lbr69 netRa69 netL69 3.016115620187341e-11
Rbbr69 netL69 node_3 -61086.300197843135
Cbr69 netL69 node_3 3.2052546359734074e-20

* Branch 70
Rabr70 node_1 netRa70 12811.992323703236
Lbr70 netRa70 netL70 2.677533072065968e-11
Rbbr70 netL70 node_3 -71420.36899549431
Cbr70 netL70 node_3 2.927905647278293e-20

* Branch 71
Rabr71 node_1 netRa71 19709.853924918156
Lbr71 netRa71 netL71 2.5543076707711532e-11
Rbbr71 netL71 node_3 -47451.61614803207
Cbr71 netL71 node_3 2.731918162797309e-20

* Branch 72
Rabr72 node_1 netRa72 16258.04306209099
Lbr72 netRa72 netL72 2.938779201214798e-11
Rbbr72 netL72 node_3 -59049.50963047863
Cbr72 netL72 node_3 3.0623020221505005e-20

* Branch 73
Rabr73 node_1 netRa73 18078.18920027984
Lbr73 netRa73 netL73 3.155388460812454e-11
Rbbr73 netL73 node_3 -58967.89648465745
Cbr73 netL73 node_3 2.9609693848549906e-20

* Branch 74
Rabr74 node_1 netRa74 21707.312989142065
Lbr74 netRa74 netL74 3.4967039989779467e-11
Rbbr74 netL74 node_3 -58465.249234754934
Cbr74 netL74 node_3 2.75590481159558e-20

* Branch 75
Rabr75 node_1 netRa75 2471.565810134102
Lbr75 netRa75 netL75 5.088629657676625e-12
Rbbr75 netL75 node_3 -15247.54361368924
Cbr75 netL75 node_3 1.3507185944198107e-19

* Branch 76
Rabr76 node_1 netRa76 -299537.2334308686
Lbr76 netRa76 netL76 2.76638979280245e-10
Rbbr76 netL76 node_3 548578.2955089498
Cbr76 netL76 node_3 1.6833086620175326e-21

* Branch 77
Rabr77 node_1 netRa77 15583.388635836392
Lbr77 netRa77 netL77 2.2156883200471633e-11
Rbbr77 netL77 node_3 -43004.34683582289
Cbr77 netL77 node_3 3.3067753812365527e-20

* Branch 78
Rabr78 node_1 netRa78 82680.68877743992
Lbr78 netRa78 netL78 8.106267233535037e-11
Rbbr78 netL78 node_3 -125706.54842274262
Cbr78 netL78 node_3 7.80015013873581e-21

* Branch 79
Rabr79 node_1 netRa79 19515.37506880497
Lbr79 netRa79 netL79 3.7411835925905326e-11
Rbbr79 netL79 node_3 -97242.47861863143
Cbr79 netL79 node_3 1.971795295914611e-20

* Branch 80
Rabr80 node_1 netRa80 26454.295899955283
Lbr80 netRa80 netL80 3.585930582883343e-11
Rbbr80 netL80 node_3 -56780.36694584179
Cbr80 netL80 node_3 2.387592418857141e-20

* Branch 81
Rabr81 node_1 netRa81 43020.218714836854
Lbr81 netRa81 netL81 4.6587410325571014e-11
Rbbr81 netL81 node_3 -71692.25710059662
Cbr81 netL81 node_3 1.5106186816852393e-20

* Branch 82
Rabr82 node_1 netRa82 35726.26393814195
Lbr82 netRa82 netL82 4.127090270190682e-11
Rbbr82 netL82 node_3 -64130.20226303533
Cbr82 netL82 node_3 1.8014335504834072e-20

* Branch 83
Rabr83 node_1 netRa83 -29465.664206628324
Lbr83 netRa83 netL83 -4.4384895175632036e-11
Rbbr83 netL83 node_3 181545.45892230235
Cbr83 netL83 node_3 -8.297280780932384e-21

* Branch 84
Rabr84 node_1 netRa84 77902.06596044956
Lbr84 netRa84 netL84 5.10062872912271e-11
Rbbr84 netL84 node_3 -93450.27301809491
Cbr84 netL84 node_3 7.006410066869863e-21

* Branch 85
Rabr85 node_1 netRa85 -228054.51624779726
Lbr85 netRa85 netL85 4.6775198938737944e-11
Rbbr85 netL85 node_3 260243.95683207596
Cbr85 netL85 node_3 7.881226200867848e-22

* Branch 86
Rabr86 node_1 netRa86 10224.078247707457
Lbr86 netRa86 netL86 2.5961718420182328e-11
Rbbr86 netL86 node_3 -84120.78830238426
Cbr86 netL86 node_3 3.0189076685117005e-20

* Branch 87
Rabr87 node_1 netRa87 10077786.600551594
Lbr87 netRa87 netL87 3.8408703213037355e-10
Rbbr87 netL87 node_3 -10085032.270937191
Cbr87 netL87 node_3 3.779096715277298e-24

* Branch 88
Rabr88 node_1 netRa88 91845.197201337
Lbr88 netRa88 netL88 2.0070939911801213e-11
Rbbr88 netL88 node_3 -104591.65109110392
Cbr88 netL88 node_3 2.0894157035050206e-21

* Branch 89
Rabr89 node_1 netRa89 4994.444863838923
Lbr89 netRa89 netL89 -1.3677925238738402e-11
Rbbr89 netL89 node_3 -21576.58047756213
Cbr89 netL89 node_3 -1.2684600496256733e-19

* Branch 90
Rabr90 node_1 netRa90 -399.30315427002546
Lbr90 netRa90 netL90 7.258545463043115e-12
Rbbr90 netL90 node_3 257480.04823439414
Cbr90 netL90 node_3 7.02759407092834e-20

* Branch 91
Rabr91 node_1 netRa91 -5320.3082479105515
Lbr91 netRa91 netL91 -1.574910191514885e-11
Rbbr91 netL91 node_3 23735.881387308134
Cbr91 netL91 node_3 -1.2480842225716895e-19

* Branch 92
Rabr92 node_1 netRa92 -527781072.8489007
Lbr92 netRa92 netL92 3.57111064054983e-09
Rbbr92 netL92 node_3 527818146.6966914
Cbr92 netL92 node_3 1.2819301955512013e-26

* Branch 93
Rabr93 node_1 netRa93 -5849547.347799878
Lbr93 netRa93 netL93 -2.273835382991589e-10
Rbbr93 netL93 node_3 5880988.783731233
Cbr93 netL93 node_3 -6.609845400286979e-24

* Branch 94
Rabr94 node_1 netRa94 -35543.001437640974
Lbr94 netRa94 netL94 2.752742221020032e-11
Rbbr94 netL94 node_3 69192.7023241725
Cbr94 netL94 node_3 1.1190195080885618e-20

* Branch 95
Rabr95 node_1 netRa95 -16939.87862755765
Lbr95 netRa95 netL95 -8.078729957014808e-12
Rbbr95 netL95 node_3 27039.277626360705
Cbr95 netL95 node_3 -1.764261150692442e-20

* Branch 96
Rabr96 node_1 netRa96 -15672.697228299521
Lbr96 netRa96 netL96 -2.965248179487541e-11
Rbbr96 netL96 node_3 85305.11796634307
Cbr96 netL96 node_3 -2.2220253464991e-20

* Branch 97
Rabr97 node_1 netRa97 -5130116.966727346
Lbr97 netRa97 netL97 -1.7011533917982827e-10
Rbbr97 netL97 node_3 5137328.034309849
Cbr97 netL97 node_3 -6.4550083658007465e-24

* Branch 98
Rabr98 node_1 netRa98 -25565.082386609338
Lbr98 netRa98 netL98 -1.1933113782979964e-11
Rbbr98 netL98 node_3 39150.17665867484
Cbr98 netL98 node_3 -1.1930138937495413e-20

* Branch 99
Rabr99 node_1 netRa99 -96673.07820432248
Lbr99 netRa99 netL99 -1.246108918235885e-11
Rbbr99 netL99 node_3 101093.72780570127
Cbr99 netL99 node_3 -1.279984468882301e-21

.ends


* Y'14
.subckt yp14 node_1 node_4
* Branch 0
Rabr0 node_1 netRa0 5654.890698947863
Lbr0 netRa0 netL0 5.610908185240118e-12
Rbbr0 netL0 node_4 -20027.446050237744
Cbr0 netL0 node_4 5.082666390364241e-20

* Branch 1
Rabr1 node_1 netRa1 -81826.98185424441
Lbr1 netRa1 netL1 -1.4595608403471468e-11
Rbbr1 netL1 node_4 89420.56226409489
Cbr1 netL1 node_4 -2.0034256901779355e-21

* Branch 2
Rabr2 node_1 netRa2 -10523.171988548793
Lbr2 netRa2 netL2 -9.842093341055195e-12
Rbbr2 netL2 node_4 29770.334602005478
Cbr2 netL2 node_4 -3.213443550108704e-20

* Branch 3
Rabr3 node_1 netRa3 -9464.121855464236
Lbr3 netRa3 netL3 -9.608001507744783e-12
Rbbr3 netL3 node_4 27530.83779262642
Cbr3 netL3 node_4 -3.776517227904172e-20

* Branch 4
Rabr4 node_1 netRa4 6750.3012174488185
Lbr4 netRa4 netL4 -9.781589336324028e-12
Rbbr4 netL4 node_4 -32414.429636891487
Cbr4 netL4 node_4 -4.3265424557906945e-20

* Branch 5
Rabr5 node_1 netRa5 2881.6595429452855
Lbr5 netRa5 netL5 -3.725362832076625e-12
Rbbr5 netL5 node_4 -17919.414019087428
Cbr5 netL5 node_4 -7.012932419741989e-20

* Branch 6
Rabr6 node_1 netRa6 7151.392521872288
Lbr6 netRa6 netL6 -5.107707731745065e-12
Rbbr6 netL6 node_4 -18185.939790418124
Cbr6 netL6 node_4 -3.866423484062914e-20

* Branch 7
Rabr7 node_1 netRa7 -26605.440662969213
Lbr7 netRa7 netL7 -8.059528547507257e-12
Rbbr7 netL7 node_4 34914.78998548567
Cbr7 netL7 node_4 -8.731388272733018e-21

* Branch 8
Rabr8 node_1 netRa8 -357376.4499615363
Lbr8 netRa8 netL8 -2.8858451631129555e-11
Rbbr8 netL8 node_4 364079.3389287274
Cbr8 netL8 node_4 -2.2216434804012553e-22

* Branch 9
Rabr9 node_1 netRa9 145812.32663766562
Lbr9 netRa9 netL9 1.7287820586672664e-11
Rbbr9 netL9 node_4 -151927.52367871604
Cbr9 netL9 node_4 7.822738570755471e-22

* Branch 10
Rabr10 node_1 netRa10 -48540.06605958189
Lbr10 netRa10 netL10 -2.1151922117737428e-11
Rbbr10 netL10 node_4 69952.6874414145
Cbr10 netL10 node_4 -6.282132963321012e-21

* Branch 11
Rabr11 node_1 netRa11 1797331.2232669431
Lbr11 netRa11 netL11 4.9619561975464865e-11
Rbbr11 netL11 node_4 -1800873.206030462
Cbr11 netL11 node_4 1.5338036396500506e-23

* Branch 12
Rabr12 node_1 netRa12 -2574.5151130346244
Lbr12 netRa12 netL12 -7.941509762560721e-12
Rbbr12 netL12 node_4 59461.819536036935
Cbr12 netL12 node_4 -5.482305435996053e-20

* Branch 13
Rabr13 node_1 netRa13 -1691.6137635700293
Lbr13 netRa13 netL13 -5.008389656887414e-12
Rbbr13 netL13 node_4 21827.376839858924
Cbr13 netL13 node_4 -1.4294373752065148e-19

* Branch 14
Rabr14 node_1 netRa14 5671.490909380743
Lbr14 netRa14 netL14 -4.8320137329065036e-12
Rbbr14 netL14 node_4 -18812.555320419182
Cbr14 netL14 node_4 -4.4640777951895863e-20

* Branch 15
Rabr15 node_1 netRa15 -54628.00270244858
Lbr15 netRa15 netL15 -1.2706373957610554e-11
Rbbr15 netL15 node_4 63224.59929290971
Cbr15 netL15 node_4 -3.692819956546524e-21

* Branch 16
Rabr16 node_1 netRa16 4003.3843029821596
Lbr16 netRa16 netL16 8.73717180755854e-12
Rbbr16 netL16 node_4 -56474.70248614423
Cbr16 netL16 node_4 4.0024923708246595e-20

* Branch 17
Rabr17 node_1 netRa17 -673719.7003706103
Lbr17 netRa17 netL17 1.455356210098557e-10
Rbbr17 netL17 node_4 691451.2554668487
Cbr17 netL17 node_4 3.1136098144433807e-22

* Branch 18
Rabr18 node_1 netRa18 1930.651654918705
Lbr18 netRa18 netL18 -3.821897720931235e-12
Rbbr18 netL18 node_4 -17749.825635435613
Cbr18 netL18 node_4 -1.0818111566971209e-19

* Branch 19
Rabr19 node_1 netRa19 647393.6724556125
Lbr19 netRa19 netL19 7.234781298372327e-11
Rbbr19 netL19 node_4 -658243.4069440282
Cbr19 netL19 node_4 1.700702983846667e-22

* Branch 20
Rabr20 node_1 netRa20 342675.31504887226
Lbr20 netRa20 netL20 -3.709161761061862e-11
Rbbr20 netL20 node_4 -351635.40166598716
Cbr20 netL20 node_4 -3.0730886570870355e-22

* Branch 21
Rabr21 node_1 netRa21 -4525.800652521131
Lbr21 netRa21 netL21 -6.6420222264227855e-12
Rbbr21 netL21 node_4 21428.671622616268
Cbr21 netL21 node_4 -7.002653266708076e-20

* Branch 22
Rabr22 node_1 netRa22 -259662.4586386414
Lbr22 netRa22 netL22 -1.7199765386614004e-11
Rbbr22 netL22 node_4 263001.58210084453
Cbr22 netL22 node_4 -2.5208225658606714e-22

* Branch 23
Rabr23 node_1 netRa23 -8244.367728158528
Lbr23 netRa23 netL23 -1.5550894142275857e-11
Rbbr23 netL23 node_4 66047.89353716308
Cbr23 netL23 node_4 -2.9235968588738494e-20

* Branch 24
Rabr24 node_1 netRa24 -43686.05291386398
Lbr24 netRa24 netL24 -2.9000111063465348e-11
Rbbr24 netL24 node_4 63698.1404193312
Cbr24 netL24 node_4 -1.0505779087110933e-20

* Branch 25
Rabr25 node_1 netRa25 -120869.12043144164
Lbr25 netRa25 netL25 -4.619274571028591e-11
Rbbr25 netL25 node_4 146397.22164598602
Cbr25 netL25 node_4 -2.6224479939433753e-21

* Branch 26
Rabr26 node_1 netRa26 221738.32379984547
Lbr26 netRa26 netL26 -6.470644633737247e-11
Rbbr26 netL26 node_4 -239064.7659907624
Cbr26 netL26 node_4 -1.216817222458843e-21

* Branch 27
Rabr27 node_1 netRa27 -59062.71960144563
Lbr27 netRa27 netL27 -3.540015052347908e-11
Rbbr27 netL27 node_4 74981.11601777129
Cbr27 netL27 node_4 -8.045092178936425e-21

* Branch 28
Rabr28 node_1 netRa28 -18382.8192927968
Lbr28 netRa28 netL28 -1.5994864740421843e-11
Rbbr28 netL28 node_4 34272.55326525573
Cbr28 netL28 node_4 -2.5615803907655358e-20

* Branch 29
Rabr29 node_1 netRa29 -9748.72355905252
Lbr29 netRa29 netL29 -1.1240520698039428e-11
Rbbr29 netL29 node_4 21213.17528960115
Cbr29 netL29 node_4 -5.496891761636677e-20

* Branch 30
Rabr30 node_1 netRa30 -42379.653761638176
Lbr30 netRa30 netL30 -2.4199485660647042e-11
Rbbr30 netL30 node_4 64230.127514311374
Cbr30 netL30 node_4 -8.93809474450415e-21

* Branch 31
Rabr31 node_1 netRa31 30552.50488280982
Lbr31 netRa31 netL31 -1.267993974680904e-11
Rbbr31 netL31 node_4 -39584.63780875074
Cbr31 netL31 node_4 -1.0444761478865038e-20

* Branch 32
Rabr32 node_1 netRa32 108010.28981499755
Lbr32 netRa32 netL32 -3.1114981887874456e-11
Rbbr32 netL32 node_4 -120187.36723194306
Cbr32 netL32 node_4 -2.3908519039743926e-21

* Branch 33
Rabr33 node_1 netRa33 -74573.81565836103
Lbr33 netRa33 netL33 -4.081463301320939e-11
Rbbr33 netL33 node_4 97002.48358679921
Cbr33 netL33 node_4 -5.669207393557278e-21

* Branch 34
Rabr34 node_1 netRa34 2184.5162864227937
Lbr34 netRa34 netL34 -5.081637460335063e-12
Rbbr34 netL34 node_4 -30304.064572115483
Cbr34 netL34 node_4 -7.524750985032102e-20

* Branch 35
Rabr35 node_1 netRa35 5702.778032174708
Lbr35 netRa35 netL35 -2.892067942929247e-12
Rbbr35 netL35 node_4 -10754.711253059742
Cbr35 netL35 node_4 -4.69503887181683e-20

* Branch 36
Rabr36 node_1 netRa36 -7869.022229445653
Lbr36 netRa36 netL36 6.1108645507086824e-12
Rbbr36 netL36 node_4 21012.758797237657
Cbr36 netL36 node_4 3.671498694299719e-20

* Branch 37
Rabr37 node_1 netRa37 -30369.59223076735
Lbr37 netRa37 netL37 -2.2950493466308106e-11
Rbbr37 netL37 node_4 44579.03895053682
Cbr37 netL37 node_4 -1.7059702796471214e-20

* Branch 38
Rabr38 node_1 netRa38 59402.63863559821
Lbr38 netRa38 netL38 -1.4189782301840202e-11
Rbbr38 netL38 node_4 -70081.3292117601
Cbr38 netL38 node_4 -3.402622037307482e-21

* Branch 39
Rabr39 node_1 netRa39 5001.041775111773
Lbr39 netRa39 netL39 -1.0079960920536635e-11
Rbbr39 netL39 node_4 -33087.636187845994
Cbr39 netL39 node_4 -6.006364156417401e-20

* Branch 40
Rabr40 node_1 netRa40 -77427.0510448541
Lbr40 netRa40 netL40 -3.267449068865053e-11
Rbbr40 netL40 node_4 98855.47151612779
Cbr40 netL40 node_4 -4.280743605428422e-21

* Branch 41
Rabr41 node_1 netRa41 33425.01783912965
Lbr41 netRa41 netL41 1.3894807063921071e-11
Rbbr41 netL41 node_4 -47522.48324258116
Cbr41 netL41 node_4 8.770938972862198e-21

* Branch 42
Rabr42 node_1 netRa42 -10576650.324134946
Lbr42 netRa42 netL42 -5.412881431464469e-10
Rbbr42 netL42 node_4 10593067.231758937
Cbr42 netL42 node_4 -4.832698896838887e-24

* Branch 43
Rabr43 node_1 netRa43 4659.999272090091
Lbr43 netRa43 netL43 -6.901884175066661e-12
Rbbr43 netL43 node_4 -26021.67658844469
Cbr43 netL43 node_4 -5.643683673407131e-20

* Branch 44
Rabr44 node_1 netRa44 -3284.589522227066
Lbr44 netRa44 netL44 -1.0938963615829456e-11
Rbbr44 netL44 node_4 47813.93768757515
Cbr44 netL44 node_4 -7.086982762807026e-20

* Branch 45
Rabr45 node_1 netRa45 125362.28600517444
Lbr45 netRa45 netL45 -2.715355175199686e-11
Rbbr45 netL45 node_4 -136883.2057731239
Cbr45 netL45 node_4 -1.5806910766769853e-21

* Branch 46
Rabr46 node_1 netRa46 -8091.096605824768
Lbr46 netRa46 netL46 9.959781782857568e-12
Rbbr46 netL46 node_4 13472.352677220842
Cbr46 netL46 node_4 9.094367125981324e-20

* Branch 47
Rabr47 node_1 netRa47 7983.759606166751
Lbr47 netRa47 netL47 -9.88759360871214e-12
Rbbr47 netL47 node_4 -25678.941228922995
Cbr47 netL47 node_4 -4.802265749036658e-20

* Branch 48
Rabr48 node_1 netRa48 19824.8119576912
Lbr48 netRa48 netL48 2.152116206925611e-11
Rbbr48 netL48 node_4 -41907.339122200516
Cbr48 netL48 node_4 2.6001552692501136e-20

* Branch 49
Rabr49 node_1 netRa49 19661.660870108415
Lbr49 netRa49 netL49 -1.610716130184904e-11
Rbbr49 netL49 node_4 -41006.04437016116
Cbr49 netL49 node_4 -1.9927347319185197e-20

* Branch 50
Rabr50 node_1 netRa50 -145894.3691341107
Lbr50 netRa50 netL50 -5.97763851318926e-11
Rbbr50 netL50 node_4 162095.51182679235
Cbr50 netL50 node_4 -2.530455074048534e-21

* Branch 51
Rabr51 node_1 netRa51 -7825.075918157371
Lbr51 netRa51 netL51 -1.3477871923777734e-11
Rbbr51 netL51 node_4 84432.13674650525
Cbr51 netL51 node_4 -2.0483815119133578e-20

* Branch 52
Rabr52 node_1 netRa52 -9727.158272695198
Lbr52 netRa52 netL52 2.4821060881593758e-11
Rbbr52 netL52 node_4 40665.53346132226
Cbr52 netL52 node_4 6.241468129450986e-20

* Branch 53
Rabr53 node_1 netRa53 3218.037554627711
Lbr53 netRa53 netL53 -8.254669214943544e-12
Rbbr53 netL53 node_4 -43543.59261991157
Cbr53 netL53 node_4 -5.861674017784178e-20

* Branch 54
Rabr54 node_1 netRa54 2515.0579000721227
Lbr54 netRa54 netL54 -1.8415018497564922e-11
Rbbr54 netL54 node_4 -156809.46094430683
Cbr54 netL54 node_4 -4.6040790334452374e-20

* Branch 55
Rabr55 node_1 netRa55 9360.758859076346
Lbr55 netRa55 netL55 -1.2952620344358224e-11
Rbbr55 netL55 node_4 -51944.05759181166
Cbr55 netL55 node_4 -2.65715949550368e-20

* Branch 56
Rabr56 node_1 netRa56 -1970.995597709734
Lbr56 netRa56 netL56 -1.299283118356651e-11
Rbbr56 netL56 node_4 108667.53720402932
Cbr56 netL56 node_4 -6.138695595411483e-20

* Branch 57
Rabr57 node_1 netRa57 482178367.1663583
Lbr57 netRa57 netL57 -1.4693738755763355e-09
Rbbr57 netL57 node_4 -482194304.09712386
Cbr57 netL57 node_4 -6.319757832648351e-27

* Branch 58
Rabr58 node_1 netRa58 4845666.978586558
Lbr58 netRa58 netL58 -2.5081826952249015e-10
Rbbr58 netL58 node_4 -4887513.785715965
Cbr58 netL58 node_4 -1.058968976987081e-23

* Branch 59
Rabr59 node_1 netRa59 155590.60330000278
Lbr59 netRa59 netL59 -6.16394929537282e-11
Rbbr59 netL59 node_4 -191968.63520907963
Cbr59 netL59 node_4 -2.0628637719439756e-21

* Branch 60
Rabr60 node_1 netRa60 -1866.1487927908427
Lbr60 netRa60 netL60 -1.5658221484828388e-11
Rbbr60 netL60 node_4 310290.6996834997
Cbr60 netL60 node_4 -2.725763596529086e-20

* Branch 61
Rabr61 node_1 netRa61 -971.5317496327738
Lbr61 netRa61 netL61 1.1767615541310376e-11
Rbbr61 netL61 node_4 74519.22469531518
Cbr61 netL61 node_4 1.6094278345567665e-19

* Branch 62
Rabr62 node_1 netRa62 -16138.941919854355
Lbr62 netRa62 netL62 -1.5035278373026185e-11
Rbbr62 netL62 node_4 39509.60613028215
Cbr62 netL62 node_4 -2.3597163688966978e-20

* Branch 63
Rabr63 node_1 netRa63 -158898.78838436044
Lbr63 netRa63 netL63 -2.8224088678948633e-11
Rbbr63 netL63 node_4 175691.04905225648
Cbr63 netL63 node_4 -1.0111366426432074e-21

* Branch 64
Rabr64 node_1 netRa64 -16472.084437098536
Lbr64 netRa64 netL64 -2.8357558110834397e-11
Rbbr64 netL64 node_4 49761.21830502807
Cbr64 netL64 node_4 -3.4629574912679013e-20

* Branch 65
Rabr65 node_1 netRa65 42840.7843908049
Lbr65 netRa65 netL65 2.2734719265488114e-11
Rbbr65 netL65 node_4 -70312.52332332154
Cbr65 netL65 node_4 7.549372018408365e-21

* Branch 66
Rabr66 node_1 netRa66 -26703.10300303148
Lbr66 netRa66 netL66 -3.668266376699972e-11
Rbbr66 netL66 node_4 62561.510861593415
Cbr66 netL66 node_4 -2.196625936179538e-20

* Branch 67
Rabr67 node_1 netRa67 -23937.332937181236
Lbr67 netRa67 netL67 -3.090382377194672e-11
Rbbr67 netL67 node_4 54798.76173688941
Cbr67 netL67 node_4 -2.3567117928179597e-20

* Branch 68
Rabr68 node_1 netRa68 -20431.270417775715
Lbr68 netRa68 netL68 -4.1756709721998924e-11
Rbbr68 netL68 node_4 106690.70780623697
Cbr68 netL68 node_4 -1.9164516391793655e-20

* Branch 69
Rabr69 node_1 netRa69 -19511.01376431713
Lbr69 netRa69 netL69 -3.0782364173827744e-11
Rbbr69 netL69 node_4 70364.66668299602
Cbr69 netL69 node_4 -2.242922709205816e-20

* Branch 70
Rabr70 node_1 netRa70 -20906.534984120273
Lbr70 netRa70 netL70 -2.3233120653852607e-11
Rbbr70 netL70 node_4 42540.33942278309
Cbr70 netL70 node_4 -2.6129293760949868e-20

* Branch 71
Rabr71 node_1 netRa71 -14598.07779113697
Lbr71 netRa71 netL71 -1.670963554348166e-11
Rbbr71 netL71 node_4 31240.745220459656
Cbr71 netL71 node_4 -3.664632605432289e-20

* Branch 72
Rabr72 node_1 netRa72 -27720.840804812666
Lbr72 netRa72 netL72 -3.0400757514109996e-11
Rbbr72 netL72 node_4 54568.14344043826
Cbr72 netL72 node_4 -2.0100763195954792e-20

* Branch 73
Rabr73 node_1 netRa73 -30466.827736861207
Lbr73 netRa73 netL73 -3.356275868563382e-11
Rbbr73 netL73 node_4 57909.34426414726
Cbr73 netL73 node_4 -1.9025798813436433e-20

* Branch 74
Rabr74 node_1 netRa74 -44656.51102851207
Lbr74 netRa74 netL74 -4.2814040949261354e-11
Rbbr74 netL74 node_4 71437.7894578529
Cbr74 netL74 node_4 -1.3421920818085491e-20

* Branch 75
Rabr75 node_1 netRa75 -260443.70339786756
Lbr75 netRa75 netL75 -7.708812768039737e-11
Rbbr75 netL75 node_4 271068.08462567476
Cbr75 netL75 node_4 -1.0919572852400685e-21

* Branch 76
Rabr76 node_1 netRa76 -47820.8918417452
Lbr76 netRa76 netL76 -4.3207996131218244e-11
Rbbr76 netL76 node_4 72175.05413143117
Cbr76 netL76 node_4 -1.25192965516847e-20

* Branch 77
Rabr77 node_1 netRa77 -30239.619196943357
Lbr77 netRa77 netL77 -2.557152966144257e-11
Rbbr77 netL77 node_4 73711.70901648572
Cbr77 netL77 node_4 -1.1472616613159445e-20

* Branch 78
Rabr78 node_1 netRa78 -66189.80916561713
Lbr78 netRa78 netL78 -4.9328294171582175e-11
Rbbr78 netL78 node_4 88089.39679804504
Cbr78 netL78 node_4 -8.460232404419691e-21

* Branch 79
Rabr79 node_1 netRa79 -241466.78980597752
Lbr79 netRa79 netL79 6.904469956943327e-11
Rbbr79 netL79 node_4 251290.87639356728
Cbr79 netL79 node_4 1.1378790014955337e-21

* Branch 80
Rabr80 node_1 netRa80 -25549.301315395245
Lbr80 netRa80 netL80 -3.685937393727053e-11
Rbbr80 netL80 node_4 83168.99297021847
Cbr80 netL80 node_4 -1.734693507795273e-20

* Branch 81
Rabr81 node_1 netRa81 -51097.75861792908
Lbr81 netRa81 netL81 -4.648379387820245e-11
Rbbr81 netL81 node_4 75127.97940834115
Cbr81 netL81 node_4 -1.2109145779363283e-20

* Branch 82
Rabr82 node_1 netRa82 159229.72437647553
Lbr82 netRa82 netL82 2.163354848456889e-10
Rbbr82 netL82 node_4 -445858.4873631082
Cbr82 netL82 node_4 3.0474816597294705e-21

* Branch 83
Rabr83 node_1 netRa83 -8451.632697396994
Lbr83 netRa83 netL83 -1.289876219961214e-11
Rbbr83 netL83 node_4 49008.62095119944
Cbr83 netL83 node_4 -3.114433636530222e-20

* Branch 84
Rabr84 node_1 netRa84 -57474.62740960144
Lbr84 netRa84 netL84 -5.74264021759597e-11
Rbbr84 netL84 node_4 88522.90006788407
Cbr84 netL84 node_4 -1.128821838663025e-20

* Branch 85
Rabr85 node_1 netRa85 -840.5149401962504
Lbr85 netRa85 netL85 -4.238236857011865e-11
Rbbr85 netL85 node_4 3795163.958166637
Cbr85 netL85 node_4 -1.3369215225107374e-20

* Branch 86
Rabr86 node_1 netRa86 -5226.321842794882
Lbr86 netRa86 netL86 -1.5818978643720762e-11
Rbbr86 netL86 node_4 58898.35011527834
Cbr86 netL86 node_4 -5.142529812234864e-20

* Branch 87
Rabr87 node_1 netRa87 1964062.6641347383
Lbr87 netRa87 netL87 -2.2479977928905893e-10
Rbbr87 netL87 node_4 -2003539.0247460199
Cbr87 netL87 node_4 -5.71254944444584e-23

* Branch 88
Rabr88 node_1 netRa88 9562.337522866079
Lbr88 netRa88 netL88 1.368167041930004e-11
Rbbr88 netL88 node_4 -17290.4741095878
Cbr88 netL88 node_4 8.278522462856708e-20

* Branch 89
Rabr89 node_1 netRa89 -2577.7493236678056
Lbr89 netRa89 netL89 7.622133020398129e-12
Rbbr89 netL89 node_4 12580.596670178455
Cbr89 netL89 node_4 2.348006816616593e-19

* Branch 90
Rabr90 node_1 netRa90 23873.7704481921
Lbr90 netRa90 netL90 -2.2384808021468236e-11
Rbbr90 netL90 node_4 -56996.63950097186
Cbr90 netL90 node_4 -1.6445266268699225e-20

* Branch 91
Rabr91 node_1 netRa91 338.05115947502736
Lbr91 netRa91 netL91 -1.1687646274726676e-11
Rbbr91 netL91 node_4 -723471.2991939598
Cbr91 netL91 node_4 -4.720901968180464e-20

* Branch 92
Rabr92 node_1 netRa92 135496.69650252222
Lbr92 netRa92 netL92 -3.403968567677997e-11
Rbbr92 netL92 node_4 -146063.48575713945
Cbr92 netL92 node_4 -1.7195830578967196e-21

* Branch 93
Rabr93 node_1 netRa93 44200.798920735084
Lbr93 netRa93 netL93 -1.754833200347113e-11
Rbbr93 netL93 node_4 -53101.556624015626
Cbr93 netL93 node_4 -7.473820684302003e-21

* Branch 94
Rabr94 node_1 netRa94 -1919.038651896004
Lbr94 netRa94 netL94 -1.006936040959021e-11
Rbbr94 netL94 node_4 149851.31549569216
Cbr94 netL94 node_4 -3.518250758031555e-20

* Branch 95
Rabr95 node_1 netRa95 8766.222921406948
Lbr95 netRa95 netL95 -1.2580576235705825e-11
Rbbr95 netL95 node_4 -60103.51907264759
Cbr95 netL95 node_4 -2.3845296990435207e-20

* Branch 96
Rabr96 node_1 netRa96 96655.42810543717
Lbr96 netRa96 netL96 1.7978322752115248e-11
Rbbr96 netL96 node_4 -105789.83656570798
Cbr96 netL96 node_4 1.7586078153214448e-21

* Branch 97
Rabr97 node_1 netRa97 103362.99305740072
Lbr97 netRa97 netL97 1.2418854686851756e-11
Rbbr97 netL97 node_4 -107360.65987918673
Cbr97 netL97 node_4 1.1193592623578344e-21

* Branch 98
Rabr98 node_1 netRa98 4997.782252118828
Lbr98 netRa98 netL98 -4.01050991070125e-12
Rbbr98 netL98 node_4 -13404.636962656541
Cbr98 netL98 node_4 -5.974432256908863e-20

* Branch 99
Rabr99 node_1 netRa99 1662.6602271295865
Lbr99 netRa99 netL99 -1.8435514962858127e-12
Rbbr99 netL99 node_4 -7567.4532014471215
Cbr99 netL99 node_4 -1.4583607976666168e-19

.ends


* Y'22
.subckt yp22 node_2 0
* Branch 0
Rabr0 node_2 netRa0 1293315.7833908445
Lbr0 netRa0 netL0 -1.6450921820165788e-10
Rbbr0 netL0 0 -1364601.568056731
Cbr0 netL0 0 -9.292069986768483e-23

* Branch 1
Rabr1 node_2 netRa1 24279.3710039378
Lbr1 netRa1 netL1 -8.702568024507145e-11
Rbbr1 netL1 0 -756832.1142179681
Cbr1 netL1 0 -4.379435700048652e-21

* Branch 2
Rabr2 node_2 netRa2 31197.695400725355
Lbr2 netRa2 netL2 -7.692425545000842e-11
Rbbr2 netL2 0 -438683.7799002283
Cbr2 netL2 0 -5.330958215894582e-21

* Branch 3
Rabr3 node_2 netRa3 275132.25777287676
Lbr3 netRa3 netL3 -7.69110180327271e-11
Rbbr3 netL3 0 -347507.0678636851
Cbr3 netL3 0 -7.995183932025439e-22

* Branch 4
Rabr4 node_2 netRa4 10761053.962443326
Lbr4 netRa4 netL4 5.765397152657606e-10
Rbbr4 netL4 0 -10842413.146975761
Cbr4 netL4 0 4.946246269786165e-24

* Branch 5
Rabr5 node_2 netRa5 67799.93719379994
Lbr5 netRa5 netL5 -2.0787861687506593e-10
Rbbr5 netL5 0 -1095368.346110444
Cbr5 netL5 0 -2.6615099489803148e-21

* Branch 6
Rabr6 node_2 netRa6 -2228.758110303673
Lbr6 netRa6 netL6 -2.0760076283348722e-10
Rbbr6 netL6 0 -53573809.527647
Cbr6 netL6 0 -4.8241574501296124e-21

* Branch 7
Rabr7 node_2 netRa7 7587.248706630143
Lbr7 netRa7 netL7 -1.4929140803821248e-10
Rbbr7 netL7 0 -2905267.2984192832
Cbr7 netL7 0 -5.323067824390763e-21

* Branch 8
Rabr8 node_2 netRa8 100073.46983679039
Lbr8 netRa8 netL8 5.613963934961518e-11
Rbbr8 netL8 0 -199020.5167122344
Cbr8 netL8 0 2.84029684850246e-21

* Branch 9
Rabr9 node_2 netRa9 -18290.399610114808
Lbr9 netRa9 netL9 -2.5073545321961654e-10
Rbbr9 netL9 0 2630925.544833956
Cbr9 netL9 0 -6.384379189329029e-21

* Branch 10
Rabr10 node_2 netRa10 4956.7626303517545
Lbr10 netRa10 netL10 -2.431385446842429e-10
Rbbr10 netL10 0 -6685218.1660743235
Cbr10 netL10 0 -4.455534397316094e-21

* Branch 11
Rabr11 node_2 netRa11 -173.39725862396787
Lbr11 netRa11 netL11 -1.7487052083010638e-10
Rbbr11 netL11 0 -17126985.670534242
Cbr11 netL11 0 -4.8344518872685156e-21

* Branch 12
Rabr12 node_2 netRa12 -8397.436065962056
Lbr12 netRa12 netL12 -1.3875076466101408e-10
Rbbr12 netL12 0 4184112.731958094
Cbr12 netL12 0 -5.014557931378853e-21

* Branch 13
Rabr13 node_2 netRa13 672903.5430992849
Lbr13 netRa13 netL13 -1.2562124832644357e-10
Rbbr13 netL13 0 -736516.6350662571
Cbr13 netL13 0 -2.5288300777129067e-22

* Branch 14
Rabr14 node_2 netRa14 139890.9391539008
Lbr14 netRa14 netL14 -5.667096754275787e-11
Rbbr14 netL14 0 -196411.07085695336
Cbr14 netL14 0 -2.0528112356592812e-21

* Branch 15
Rabr15 node_2 netRa15 20055.62744579073
Lbr15 netRa15 netL15 -2.2964308482282165e-10
Rbbr15 netL15 0 -1318543.591283623
Cbr15 netL15 0 -7.713882035731241e-21

* Branch 16
Rabr16 node_2 netRa16 17487.456911033143
Lbr16 netRa16 netL16 -1.3105881768758062e-10
Rbbr16 netL16 0 -1783959.9675902468
Cbr16 netL16 0 -3.888024249553592e-21

* Branch 17
Rabr17 node_2 netRa17 483922.31475869217
Lbr17 netRa17 netL17 1.0483903434023538e-10
Rbbr17 netL17 0 -549445.7592113393
Cbr17 netL17 0 3.9515827995304014e-22

* Branch 18
Rabr18 node_2 netRa18 62511.737020271066
Lbr18 netRa18 netL18 -2.9458516827685194e-10
Rbbr18 netL18 0 -990168.4467354722
Cbr18 netL18 0 -4.553138054915818e-21

* Branch 19
Rabr19 node_2 netRa19 103134.55896391647
Lbr19 netRa19 netL19 5.24659401525772e-11
Rbbr19 netL19 0 -195083.31082428043
Cbr19 netL19 0 2.620253228938087e-21

* Branch 20
Rabr20 node_2 netRa20 -183438.7038556616
Lbr20 netRa20 netL20 -2.979121932171733e-10
Rbbr20 netL20 0 866058.571054558
Cbr20 netL20 0 -1.9014721806338568e-21

* Branch 21
Rabr21 node_2 netRa21 44070.79485124663
Lbr21 netRa21 netL21 -1.0001859929869583e-10
Rbbr21 netL21 0 -671811.6966477963
Cbr21 netL21 0 -3.31581554646152e-21

* Branch 22
Rabr22 node_2 netRa22 2532.7325143518574
Lbr22 netRa22 netL22 -1.859351047096071e-10
Rbbr22 netL22 0 -9372851.360132517
Cbr22 netL22 0 -4.986323180530441e-21

* Branch 23
Rabr23 node_2 netRa23 102352.60880342383
Lbr23 netRa23 netL23 -2.3653513345274386e-10
Rbbr23 netL23 0 -367092.8554007521
Cbr23 netL23 0 -6.190145456073788e-21

* Branch 24
Rabr24 node_2 netRa24 32266.859477655176
Lbr24 netRa24 netL24 -3.709972565815412e-11
Rbbr24 netL24 0 -159370.56862415757
Cbr24 netL24 0 -7.155374945355562e-21

* Branch 25
Rabr25 node_2 netRa25 2330041418.9551377
Lbr25 netRa25 netL25 -7.745833547118339e-09
Rbbr25 netL25 0 -2330120822.8470154
Cbr25 netL25 0 -1.4266452186307534e-27

* Branch 26
Rabr26 node_2 netRa26 -342911.6778873737
Lbr26 netRa26 netL26 -3.3455934433991107e-10
Rbbr26 netL26 0 837440.0794215943
Cbr26 netL26 0 -1.1727888868129377e-21

* Branch 27
Rabr27 node_2 netRa27 -18942.723472516966
Lbr27 netRa27 netL27 -1.7029267452683158e-10
Rbbr27 netL27 0 1359668.7221562609
Cbr27 netL27 0 -7.034140066702328e-21

* Branch 28
Rabr28 node_2 netRa28 -27414.56379768869
Lbr28 netRa28 netL28 -2.563293415185485e-10
Rbbr28 netL28 0 1947497.7503188164
Cbr28 netL28 0 -5.084838553545676e-21

* Branch 29
Rabr29 node_2 netRa29 1113519.5680085998
Lbr29 netRa29 netL29 -2.1887056791652477e-10
Rbbr29 netL29 0 -1181761.7945340986
Cbr29 netL29 0 -1.661320914334767e-22

* Branch 30
Rabr30 node_2 netRa30 -90095346.38694057
Lbr30 netRa30 netL30 5.601439561004875e-09
Rbbr30 netL30 0 91225215.14892055
Cbr30 netL30 0 6.812758996525962e-25

* Branch 31
Rabr31 node_2 netRa31 -688236.5597125662
Lbr31 netRa31 netL31 -3.8212643173297236e-10
Rbbr31 netL31 0 1382279.3695070993
Cbr31 netL31 0 -4.029695774386457e-22

* Branch 32
Rabr32 node_2 netRa32 94456127.16203412
Lbr32 netRa32 netL32 2.122880473677471e-09
Rbbr32 netL32 0 -94521048.68807422
Cbr32 netL32 0 2.378050685839763e-25

* Branch 33
Rabr33 node_2 netRa33 -22608.231282571323
Lbr33 netRa33 netL33 -2.326423911391434e-11
Rbbr33 netL33 0 105886.06676975173
Cbr33 netL33 0 -9.771327257122884e-21

* Branch 34
Rabr34 node_2 netRa34 113265.83078336637
Lbr34 netRa34 netL34 -7.091157402509362e-11
Rbbr34 netL34 0 -221176.22698806337
Cbr34 netL34 0 -2.8220861386507785e-21

* Branch 35
Rabr35 node_2 netRa35 -2339.637027149434
Lbr35 netRa35 netL35 -4.784630447821567e-11
Rbbr35 netL35 0 3208080.680220392
Cbr35 netL35 0 -7.051571239808414e-21

* Branch 36
Rabr36 node_2 netRa36 -220252.09557167592
Lbr36 netRa36 netL36 -2.1129239600519574e-10
Rbbr36 netL36 0 527603.1983995435
Cbr36 netL36 0 -1.8259136285552362e-21

* Branch 37
Rabr37 node_2 netRa37 24245.826636461465
Lbr37 netRa37 netL37 -4.664433963579909e-11
Rbbr37 netL37 0 -237660.3866540446
Cbr37 netL37 0 -8.031559117576683e-21

* Branch 38
Rabr38 node_2 netRa38 285550.30247347074
Lbr38 netRa38 netL38 -2.353404796107937e-10
Rbbr38 netL38 0 -411619.8175469563
Cbr38 netL38 0 -1.996122267928428e-21

* Branch 39
Rabr39 node_2 netRa39 1238129.7700038764
Lbr39 netRa39 netL39 4.760966280231603e-10
Rbbr39 netL39 0 -1347369.361306162
Cbr39 netL39 0 2.8577938549224646e-22

* Branch 40
Rabr40 node_2 netRa40 51815.762507110674
Lbr40 netRa40 netL40 -1.1726485024051565e-10
Rbbr40 netL40 0 -231253.39294832613
Cbr40 netL40 0 -9.712227969013758e-21

* Branch 41
Rabr41 node_2 netRa41 93793.01527675119
Lbr41 netRa41 netL41 -1.2544841888586326e-10
Rbbr41 netL41 0 -233907.1341227181
Cbr41 netL41 0 -5.6927989644523374e-21

* Branch 42
Rabr42 node_2 netRa42 -10225.38662534709
Lbr42 netRa42 netL42 -1.0823195110822313e-10
Rbbr42 netL42 0 2465477.585749482
Cbr42 netL42 0 -4.4150219216833665e-21

* Branch 43
Rabr43 node_2 netRa43 21838.869404375753
Lbr43 netRa43 netL43 -5.93807961357585e-11
Rbbr43 netL43 0 -267474.1992660631
Cbr43 netL43 0 -1.0096219852755505e-20

* Branch 44
Rabr44 node_2 netRa44 57573.09364541691
Lbr44 netRa44 netL44 -1.1068936985338706e-10
Rbbr44 netL44 0 -461869.18860361463
Cbr44 netL44 0 -4.1450691290223815e-21

* Branch 45
Rabr45 node_2 netRa45 -83543381.89868215
Lbr45 netRa45 netL45 1.1318415384178528e-09
Rbbr45 netL45 0 83585643.23215035
Cbr45 netL45 0 1.6207998980277352e-25

* Branch 46
Rabr46 node_2 netRa46 206664.15969234877
Lbr46 netRa46 netL46 -1.9251652475601103e-10
Rbbr46 netL46 0 -362755.72644718096
Cbr46 netL46 0 -2.562973540723886e-21

* Branch 47
Rabr47 node_2 netRa47 76990.84584863149
Lbr47 netRa47 netL47 -9.599470642490328e-11
Rbbr47 netL47 0 -335919.29648063803
Cbr47 netL47 0 -3.702759662216555e-21

* Branch 48
Rabr48 node_2 netRa48 206446.22871178557
Lbr48 netRa48 netL48 -2.108941620932665e-10
Rbbr48 netL48 0 -447804.73126232263
Cbr48 netL48 0 -2.277243369191241e-21

* Branch 49
Rabr49 node_2 netRa49 -35379.027373776866
Lbr49 netRa49 netL49 -7.209655166507643e-11
Rbbr49 netL49 0 519902.09053061315
Cbr49 netL49 0 -3.93327119783393e-21

* Branch 50
Rabr50 node_2 netRa50 4732.706916924267
Lbr50 netRa50 netL50 -1.4648224734535732e-10
Rbbr50 netL50 0 -7901357.998851566
Cbr50 netL50 0 -3.722951110646914e-21

* Branch 51
Rabr51 node_2 netRa51 229324.49427290214
Lbr51 netRa51 netL51 -1.7375307896016016e-10
Rbbr51 netL51 0 -419677.93629019987
Cbr51 netL51 0 -1.803501539303483e-21

* Branch 52
Rabr52 node_2 netRa52 22811.61245737456
Lbr52 netRa52 netL52 -1.039058878256374e-10
Rbbr52 netL52 0 -1017431.4417488754
Cbr52 netL52 0 -4.449607623073035e-21

* Branch 53
Rabr53 node_2 netRa53 121694.88171243115
Lbr53 netRa53 netL53 -2.360607095267304e-10
Rbbr53 netL53 0 -356970.3859572855
Cbr53 netL53 0 -5.421169488002858e-21

* Branch 54
Rabr54 node_2 netRa54 75759.02006074558
Lbr54 netRa54 netL54 -2.124312049190393e-10
Rbbr54 netL54 0 -719506.8940766371
Cbr54 netL54 0 -3.884525066740796e-21

* Branch 55
Rabr55 node_2 netRa55 299434.4146910186
Lbr55 netRa55 netL55 3.2594023693320715e-10
Rbbr55 netL55 0 -552582.6519049441
Cbr55 netL55 0 1.9723467265199235e-21

* Branch 56
Rabr56 node_2 netRa56 320979.15928780433
Lbr56 netRa56 netL56 -2.472592283790359e-10
Rbbr56 netL56 0 -571886.7339864178
Cbr56 netL56 0 -1.3460495349072298e-21

* Branch 57
Rabr57 node_2 netRa57 21251.969528037822
Lbr57 netRa57 netL57 -2.1966255557708677e-10
Rbbr57 netL57 0 -1067903.3883378704
Cbr57 netL57 0 -9.596043513892407e-21

* Branch 58
Rabr58 node_2 netRa58 456743.4513344639
Lbr58 netRa58 netL58 -3.8237267124642676e-10
Rbbr58 netL58 0 -746241.0485117608
Cbr58 netL58 0 -1.1210794280701856e-21

* Branch 59
Rabr59 node_2 netRa59 -92190.21702212583
Lbr59 netRa59 netL59 1.6818643336433058e-10
Rbbr59 netL59 0 910075.5590392848
Cbr59 netL59 0 2.0016811783939084e-21

* Branch 60
Rabr60 node_2 netRa60 160556.9884544901
Lbr60 netRa60 netL60 9.383310460275489e-11
Rbbr60 netL60 0 -355907.013312046
Cbr60 netL60 0 1.6427654682041626e-21

* Branch 61
Rabr61 node_2 netRa61 48191.13896625609
Lbr61 netRa61 netL61 -1.4703893971307485e-10
Rbbr61 netL61 0 -621039.4516130624
Cbr61 netL61 0 -4.9041904091687266e-21

* Branch 62
Rabr62 node_2 netRa62 1812936.6516713712
Lbr62 netRa62 netL62 7.236190939483122e-10
Rbbr62 netL62 0 -2653037.9385027005
Cbr62 netL62 0 1.5048077130597139e-22

* Branch 63
Rabr63 node_2 netRa63 559291.3606529493
Lbr63 netRa63 netL63 -5.011360473557368e-10
Rbbr63 netL63 0 -814097.5443396907
Cbr63 netL63 0 -1.1000786140751971e-21

* Branch 64
Rabr64 node_2 netRa64 887827276.5541828
Lbr64 netRa64 netL64 9.780632922752796e-09
Rbbr64 netL64 0 -888002216.9692227
Cbr64 netL64 0 1.2405864637578724e-26

* Branch 65
Rabr65 node_2 netRa65 53576.17952059391
Lbr65 netRa65 netL65 -1.7059525986904223e-10
Rbbr65 netL65 0 -1144289.1892947832
Cbr65 netL65 0 -2.7780966308416494e-21

* Branch 66
Rabr66 node_2 netRa66 -19812.578562863317
Lbr66 netRa66 netL66 -1.1054156011757293e-10
Rbbr66 netL66 0 1306234.0019042778
Cbr66 netL66 0 -4.283608149254295e-21

* Branch 67
Rabr67 node_2 netRa67 36309.77780954985
Lbr67 netRa67 netL67 -2.752834406395526e-10
Rbbr67 netL67 0 -904111.4257978336
Cbr67 netL67 0 -8.358422955635161e-21

* Branch 68
Rabr68 node_2 netRa68 25262.97643152702
Lbr68 netRa68 netL68 -1.8578135894218888e-10
Rbbr68 netL68 0 -2560720.3861846263
Cbr68 netL68 0 -2.863097092866114e-21

* Branch 69
Rabr69 node_2 netRa69 -234461.3355511518
Lbr69 netRa69 netL69 1.3359184973609262e-10
Rbbr69 netL69 0 475155.5776325305
Cbr69 netL69 0 1.1988868075465308e-21

* Branch 70
Rabr70 node_2 netRa70 43463.29488448357
Lbr70 netRa70 netL70 -2.2777238866281557e-10
Rbbr70 netL70 0 -688025.8163851176
Cbr70 netL70 0 -7.602916140153738e-21

* Branch 71
Rabr71 node_2 netRa71 109325.34939116707
Lbr71 netRa71 netL71 -3.2428552168605726e-10
Rbbr71 netL71 0 -1299580.9006619176
Cbr71 netL71 0 -2.2805863001757544e-21

* Branch 72
Rabr72 node_2 netRa72 181680.44159158316
Lbr72 netRa72 netL72 -4.212834388505673e-10
Rbbr72 netL72 0 -1812802.3004213755
Cbr72 netL72 0 -1.2783183564250369e-21

* Branch 73
Rabr73 node_2 netRa73 88831.11742271109
Lbr73 netRa73 netL73 -3.279668924086401e-10
Rbbr73 netL73 0 -2166873.216580628
Cbr73 netL73 0 -1.702561765065399e-21

* Branch 74
Rabr74 node_2 netRa74 -12461.346057116123
Lbr74 netRa74 netL74 -9.416965614894768e-11
Rbbr74 netL74 0 359921.3345984536
Cbr74 netL74 0 -2.1005953750921622e-20

* Branch 75
Rabr75 node_2 netRa75 120122.77567685404
Lbr75 netRa75 netL75 -5.365012809762105e-10
Rbbr75 netL75 0 -2371065.1589065366
Cbr75 netL75 0 -1.883443306139895e-21

* Branch 76
Rabr76 node_2 netRa76 -27976.577297184172
Lbr76 netRa76 netL76 -3.6649400830966817e-10
Rbbr76 netL76 0 2144617.591587868
Cbr76 netL76 0 -6.109528461532046e-21

* Branch 77
Rabr77 node_2 netRa77 -18128.798236939834
Lbr77 netRa77 netL77 -2.826855200389569e-10
Rbbr77 netL77 0 1758414.7262006595
Cbr77 netL77 0 -8.868072535535846e-21

* Branch 78
Rabr78 node_2 netRa78 -749008.2110683267
Lbr78 netRa78 netL78 -6.434906259168455e-10
Rbbr78 netL78 0 1524929.9999261089
Cbr78 netL78 0 -5.633894309733342e-22

* Branch 79
Rabr79 node_2 netRa79 28750.361904212747
Lbr79 netRa79 netL79 -8.253447881153731e-10
Rbbr79 netL79 0 -19090598.166173182
Cbr79 netL79 0 -1.5019725160088683e-21

* Branch 80
Rabr80 node_2 netRa80 234165.72751221966
Lbr80 netRa80 netL80 -5.993821204677889e-10
Rbbr80 netL80 0 -1729239.1210393498
Cbr80 netL80 0 -1.4799984062352537e-21

* Branch 81
Rabr81 node_2 netRa81 181123.6479846241
Lbr81 netRa81 netL81 -7.056745810912452e-10
Rbbr81 netL81 0 -2307289.6065528663
Cbr81 netL81 0 -1.6881278253962518e-21

* Branch 82
Rabr82 node_2 netRa82 286474.3523018379
Lbr82 netRa82 netL82 -4.610470290985148e-10
Rbbr82 netL82 0 -1175843.2634381815
Cbr82 netL82 0 -1.3684535713987634e-21

* Branch 83
Rabr83 node_2 netRa83 85742002.24423714
Lbr83 netRa83 netL83 -1.203947677011852e-08
Rbbr83 netL83 0 -86997208.24517865
Cbr83 netL83 0 -1.6139929856757049e-24

* Branch 84
Rabr84 node_2 netRa84 1128946.8007025952
Lbr84 netRa84 netL84 -9.39027854661205e-10
Rbbr84 netL84 0 -2034869.568896753
Cbr84 netL84 0 -4.087158235693788e-22

* Branch 85
Rabr85 node_2 netRa85 -350707.85645228
Lbr85 netRa85 netL85 1.4311158904733716e-10
Rbbr85 netL85 0 487036.9568122854
Cbr85 netL85 0 8.378041026585834e-22

* Branch 86
Rabr86 node_2 netRa86 3686244.470982048
Lbr86 netRa86 netL86 -2.2638006539884653e-09
Rbbr86 netL86 0 -4553401.613515008
Cbr86 netL86 0 -1.3485743985416287e-22

* Branch 87
Rabr87 node_2 netRa87 2396097.76416512
Lbr87 netRa87 netL87 8.46691276798524e-10
Rbbr87 netL87 0 -2924112.4421717566
Cbr87 netL87 0 1.208523102505619e-22

* Branch 88
Rabr88 node_2 netRa88 5785271.375219854
Lbr88 netRa88 netL88 -1.7382205383021485e-09
Rbbr88 netL88 0 -6312971.29652857
Cbr88 netL88 0 -4.7590792172141124e-23

* Branch 89
Rabr89 node_2 netRa89 -58249.41088229939
Lbr89 netRa89 netL89 -7.725000464736028e-11
Rbbr89 netL89 0 302024.4294283789
Cbr89 netL89 0 -4.3922473395606864e-21

* Branch 90
Rabr90 node_2 netRa90 -190304.72892763957
Lbr90 netRa90 netL90 4.808370509858991e-10
Rbbr90 netL90 0 1462269.125703686
Cbr90 netL90 0 1.7269356563292972e-21

* Branch 91
Rabr91 node_2 netRa91 -72412.04386103961
Lbr91 netRa91 netL91 2.9641905295544876e-10
Rbbr91 netL91 0 2270063.0890721795
Cbr91 netL91 0 1.8014441148247178e-21

* Branch 92
Rabr92 node_2 netRa92 -54187.8651811539
Lbr92 netRa92 netL92 1.1678473746880707e-10
Rbbr92 netL92 0 865740.5713467859
Cbr92 netL92 0 2.487880862050543e-21

* Branch 93
Rabr93 node_2 netRa93 -368999.9364941958
Lbr93 netRa93 netL93 3.2718673184407846e-10
Rbbr93 netL93 0 937788.0016947265
Cbr93 netL93 0 9.452105432879139e-22

* Branch 94
Rabr94 node_2 netRa94 -623513.2423806184
Lbr94 netRa94 netL94 2.9903239432759757e-10
Rbbr94 netL94 0 941955.8562522125
Cbr94 netL94 0 5.090077056941226e-22

* Branch 95
Rabr95 node_2 netRa95 -100394.72470117349
Lbr95 netRa95 netL95 1.2752246370429114e-10
Rbbr95 netL95 0 434423.2296009227
Cbr95 netL95 0 2.9212296161762283e-21

* Branch 96
Rabr96 node_2 netRa96 -308977.9000565247
Lbr96 netRa96 netL96 1.6397807687099142e-10
Rbbr96 netL96 0 506872.9276195187
Cbr96 netL96 0 1.0466120887628396e-21

* Branch 97
Rabr97 node_2 netRa97 -223427.84499719567
Lbr97 netRa97 netL97 1.2979077046658822e-10
Rbbr97 netL97 0 416205.773528606
Cbr97 netL97 0 1.3950775881313893e-21

* Branch 98
Rabr98 node_2 netRa98 -18923.080121584746
Lbr98 netRa98 netL98 4.650147485714509e-11
Rbbr98 netL98 0 189159.60537923622
Cbr98 netL98 0 1.2959305412201474e-20

* Branch 99
Rabr99 node_2 netRa99 -171691071.95114645
Lbr99 netRa99 netL99 1.6525242320865315e-09
Rbbr99 netL99 0 171734909.3164085
Cbr99 netL99 0 5.604422410004575e-26

.ends


* Y'23
.subckt yp23 node_2 node_3
* Branch 0
Rabr0 node_2 netRa0 -1738788.060093933
Lbr0 netRa0 netL0 -7.118808035712333e-11
Rbbr0 netL0 node_3 1747255.5236566078
Cbr0 netL0 node_3 -2.345602392157779e-23

* Branch 1
Rabr1 node_2 netRa1 1963.0497319894166
Lbr1 netRa1 netL1 5.361173263435794e-12
Rbbr1 netL1 node_3 -41409.24394546155
Cbr1 netL1 node_3 7.060189290221652e-20

* Branch 2
Rabr2 node_2 netRa2 -12922.411662417846
Lbr2 netRa2 netL2 -1.101206773211705e-11
Rbbr2 netL2 node_3 30280.02874166599
Cbr2 netL2 node_3 -2.8711901446929526e-20

* Branch 3
Rabr3 node_2 netRa3 11568.506296002372
Lbr3 netRa3 netL3 -1.127396727833347e-11
Rbbr3 netL3 node_3 -31730.040501853662
Cbr3 netL3 node_3 -3.005205708857534e-20

* Branch 4
Rabr4 node_2 netRa4 582.6101358305895
Lbr4 netRa4 netL4 -2.8127230448871384e-12
Rbbr4 netL4 node_3 -39850.32207060647
Cbr4 netL4 node_3 -1.0926427809181593e-19

* Branch 5
Rabr5 node_2 netRa5 -22576.405225039976
Lbr5 netRa5 netL5 -1.526051350052556e-11
Rbbr5 netL5 node_3 44015.66888137882
Cbr5 netL5 node_3 -1.5592941520887655e-20

* Branch 6
Rabr6 node_2 netRa6 -769456.4494416305
Lbr6 netRa6 netL6 -4.5048584776148925e-11
Rbbr6 netL6 node_3 777058.7516065935
Cbr6 netL6 node_3 -7.544092706067161e-23

* Branch 7
Rabr7 node_2 netRa7 2832.6556729566146
Lbr7 netRa7 netL7 -3.8614417068673766e-12
Rbbr7 netL7 node_3 -18495.661591107924
Cbr7 netL7 node_3 -7.158088339918248e-20

* Branch 8
Rabr8 node_2 netRa8 -233920.35081980718
Lbr8 netRa8 netL8 2.1882655077929982e-11
Rbbr8 netL8 node_3 239889.4927662748
Cbr8 netL8 node_3 3.893175904938461e-22

* Branch 9
Rabr9 node_2 netRa9 -28835.704439788533
Lbr9 netRa9 netL9 -8.062519104429269e-12
Rbbr9 netL9 node_3 36514.163211519895
Cbr9 netL9 node_3 -7.694802294825361e-21

* Branch 10
Rabr10 node_2 netRa10 -2879.577573798832
Lbr10 netRa10 netL10 -6.5772988508534085e-12
Rbbr10 netL10 node_3 23056.35154015646
Cbr10 netL10 node_3 -1.0313841015097288e-19

* Branch 11
Rabr11 node_2 netRa11 100143.6921603974
Lbr11 netRa11 netL11 1.2517468217022626e-11
Rbbr11 netL11 node_3 -104193.62524624109
Cbr11 netL11 node_3 1.2021973874209457e-21

* Branch 12
Rabr12 node_2 netRa12 7586.148592653121
Lbr12 netRa12 netL12 -3.9647445083216225e-12
Rbbr12 netL12 node_3 -13678.055325107112
Cbr12 netL12 node_3 -3.7874529730762783e-20

* Branch 13
Rabr13 node_2 netRa13 -147220.83316240436
Lbr13 netRa13 netL13 -2.2703775722905657e-11
Rbbr13 netL13 node_3 157385.4284006427
Cbr13 netL13 node_3 -9.823554196798536e-22

* Branch 14
Rabr14 node_2 netRa14 -2447.640109972564
Lbr14 netRa14 netL14 -7.579794723266793e-12
Rbbr14 netL14 node_3 56860.447297759965
Cbr14 netL14 node_3 -5.737047778762177e-20

* Branch 15
Rabr15 node_2 netRa15 -340781.51563186984
Lbr15 netRa15 netL15 -6.343912231598717e-11
Rbbr15 netL15 node_3 368075.217572289
Cbr15 netL15 node_3 -5.072878426313439e-22

* Branch 16
Rabr16 node_2 netRa16 2092.2333942088762
Lbr16 netRa16 netL16 5.5650791878606724e-12
Rbbr16 netL16 node_3 -42870.08768686712
Cbr16 netL16 node_3 6.448625976056349e-20

* Branch 17
Rabr17 node_2 netRa17 204764.3028037766
Lbr17 netRa17 netL17 -4.8928742065182844e-11
Rbbr17 netL17 node_3 -220379.7513776247
Cbr17 netL17 node_3 -1.080745655318618e-21

* Branch 18
Rabr18 node_2 netRa18 -760520.4893793251
Lbr18 netRa18 netL18 -1.4284593198189592e-10
Rbbr18 netL18 node_3 799226.78560737
Cbr18 netL18 node_3 -2.355974903285498e-22

* Branch 19
Rabr19 node_2 netRa19 -18329.058658958376
Lbr19 netRa19 netL19 -3.128169411196714e-11
Rbbr19 netL19 node_3 123745.97787599756
Cbr19 netL19 node_3 -1.4104177377774617e-20

* Branch 20
Rabr20 node_2 netRa20 2422.5886330867966
Lbr20 netRa20 netL20 -4.230438594892199e-12
Rbbr20 netL20 node_3 -18024.36030434532
Cbr20 netL20 node_3 -9.478075353998585e-20

* Branch 21
Rabr21 node_2 netRa21 -28018.449272102287
Lbr21 netRa21 netL21 -1.958388050382119e-11
Rbbr21 netL21 node_3 43792.16727157432
Cbr21 netL21 node_3 -1.6102127306439525e-20

* Branch 22
Rabr22 node_2 netRa22 -4265.640472288468
Lbr22 netRa22 netL22 -6.392012058025727e-12
Rbbr22 netL22 node_3 20900.033718719606
Cbr22 netL22 node_3 -7.305711247989386e-20

* Branch 23
Rabr23 node_2 netRa23 -41799.37854564811
Lbr23 netRa23 netL23 -2.3963992363030686e-11
Rbbr23 netL23 node_3 63650.902767558495
Cbr23 netL23 node_3 -9.068914199294627e-21

* Branch 24
Rabr24 node_2 netRa24 -2287620.7956419894
Lbr24 netRa24 netL24 -2.718200808185032e-10
Rbbr24 netL24 node_3 2305880.9094901807
Cbr24 netL24 node_3 -5.1602825727774407e-23

* Branch 25
Rabr25 node_2 netRa25 84154086.41294718
Lbr25 netRa25 netL25 -5.262617230061417e-10
Rbbr25 netL25 node_3 -84161442.92254964
Cbr25 netL25 node_3 -7.429869641969551e-26

* Branch 26
Rabr26 node_2 netRa26 -27677.894252615602
Lbr26 netRa26 netL26 -1.879735465676052e-11
Rbbr26 netL26 node_3 38945.15530852918
Cbr26 netL26 node_3 -1.7578345399149588e-20

* Branch 27
Rabr27 node_2 netRa27 3863.3275935700194
Lbr27 netRa27 netL27 -4.173166247345497e-12
Rbbr27 netL27 node_3 -18358.91794240694
Cbr27 netL27 node_3 -5.810690767657578e-20

* Branch 28
Rabr28 node_2 netRa28 138377.37125457253
Lbr28 netRa28 netL28 -3.562463442855141e-11
Rbbr28 netL28 node_3 -150833.36799540304
Cbr28 netL28 node_3 -1.7019452070992792e-21

* Branch 29
Rabr29 node_2 netRa29 -1179.151829832826
Lbr29 netRa29 netL29 -4.229830254889674e-12
Rbbr29 netL29 node_3 39353.5133617214
Cbr29 netL29 node_3 -9.488408032586213e-20

* Branch 30
Rabr30 node_2 netRa30 -131207.7603629776
Lbr30 netRa30 netL30 -5.539638583413619e-11
Rbbr30 netL30 node_3 148726.05486940435
Cbr30 netL30 node_3 -2.8517908003074575e-21

* Branch 31
Rabr31 node_2 netRa31 -80216.78012841631
Lbr31 netRa31 netL31 -3.937454166773513e-11
Rbbr31 netL31 node_3 100457.1770481099
Cbr31 netL31 node_3 -4.91208320238263e-21

* Branch 32
Rabr32 node_2 netRa32 -118621.10676463686
Lbr32 netRa32 netL32 -4.149917202445545e-11
Rbbr32 netL32 node_3 141144.30435988508
Cbr32 netL32 node_3 -2.486969931862297e-21

* Branch 33
Rabr33 node_2 netRa33 18884.639557562037
Lbr33 netRa33 netL33 -1.1269821614699939e-11
Rbbr33 netL33 node_3 -30416.561447366275
Cbr33 netL33 node_3 -1.951377348923652e-20

* Branch 34
Rabr34 node_2 netRa34 17558.544770025517
Lbr34 netRa34 netL34 -1.7920858698640987e-11
Rbbr34 netL34 node_3 -34203.767018957966
Cbr34 netL34 node_3 -2.956890387884535e-20

* Branch 35
Rabr35 node_2 netRa35 18164.20787791067
Lbr35 netRa35 netL35 -7.426498417089749e-12
Rbbr35 netL35 node_3 -27700.634606231597
Cbr35 netL35 node_3 -1.4707467031874227e-20

* Branch 36
Rabr36 node_2 netRa36 -153376.81549756727
Lbr36 netRa36 netL36 -5.955734859237455e-11
Rbbr36 netL36 node_3 176465.80974765363
Cbr36 netL36 node_3 -2.2075697837656774e-21

* Branch 37
Rabr37 node_2 netRa37 -85658.32479801512
Lbr37 netRa37 netL37 -4.006400394501593e-11
Rbbr37 netL37 node_3 100961.14574453025
Cbr37 netL37 node_3 -4.6504792090444575e-21

* Branch 38
Rabr38 node_2 netRa38 6940.0841571875135
Lbr38 netRa38 netL38 -3.339593356373833e-12
Rbbr38 netL38 node_3 -12479.053928451509
Cbr38 netL38 node_3 -3.8410495875047146e-20

* Branch 39
Rabr39 node_2 netRa39 -10922.90310661292
Lbr39 netRa39 netL39 6.217169208431655e-12
Rbbr39 netL39 node_3 20751.332836716414
Cbr39 netL39 node_3 2.730421504117849e-20

* Branch 40
Rabr40 node_2 netRa40 -494164.4349847831
Lbr40 netRa40 netL40 -1.2255943956333229e-10
Rbbr40 netL40 node_3 512331.4263556941
Cbr40 netL40 node_3 -4.849988004888776e-22

* Branch 41
Rabr41 node_2 netRa41 2840.333865337993
Lbr41 netRa41 netL41 -1.080097921725972e-11
Rbbr41 netL41 node_3 -58881.68956876685
Cbr41 netL41 node_3 -6.286108274940825e-20

* Branch 42
Rabr42 node_2 netRa42 171955.0224874705
Lbr42 netRa42 netL42 -3.658061912397028e-11
Rbbr42 netL42 node_3 -184580.95883111292
Cbr42 netL42 node_3 -1.151092720752987e-21

* Branch 43
Rabr43 node_2 netRa43 19652.56249822478
Lbr43 netRa43 netL43 2.529493325569637e-11
Rbbr43 netL43 node_3 -50541.84498063808
Cbr43 netL43 node_3 2.5651902649207567e-20

* Branch 44
Rabr44 node_2 netRa44 -95921.2399568918
Lbr44 netRa44 netL44 4.499045701297595e-11
Rbbr44 netL44 node_3 105182.81788935317
Cbr44 netL44 node_3 4.448248614231311e-21

* Branch 45
Rabr45 node_2 netRa45 22852.893697790532
Lbr45 netRa45 netL45 1.4736165429481407e-11
Rbbr45 netL45 node_3 -46102.706529632625
Cbr45 netL45 node_3 1.4032230971904072e-20

* Branch 46
Rabr46 node_2 netRa46 -33694.56173873887
Lbr46 netRa46 netL46 4.604433948777642e-11
Rbbr46 netL46 node_3 64324.257395791974
Cbr46 netL46 node_3 2.1110062258910532e-20

* Branch 47
Rabr47 node_2 netRa47 -2690.029503352507
Lbr47 netRa47 netL47 3.188270384068457e-11
Rbbr47 netL47 node_3 189281.64373955937
Cbr47 netL47 node_3 5.939488805615976e-20

* Branch 48
Rabr48 node_2 netRa48 3489.4375675717315
Lbr48 netRa48 netL48 -7.664348270559654e-12
Rbbr48 netL48 node_3 -38661.40807622484
Cbr48 netL48 node_3 -5.62846592621201e-20

* Branch 49
Rabr49 node_2 netRa49 494751.78881903604
Lbr49 netRa49 netL49 -5.658016818501162e-11
Rbbr49 netL49 node_3 -507440.7729115335
Cbr49 netL49 node_3 -2.2526537178237076e-22

* Branch 50
Rabr50 node_2 netRa50 -1069.8710524165267
Lbr50 netRa50 netL50 -8.410138721117909e-12
Rbbr50 netL50 node_3 82873.17141748701
Cbr50 netL50 node_3 -9.766879501882175e-20

* Branch 51
Rabr51 node_2 netRa51 6547.395021971895
Lbr51 netRa51 netL51 -1.1073382629883088e-11
Rbbr51 netL51 node_3 -33580.63377088157
Cbr51 netL51 node_3 -5.013114724461992e-20

* Branch 52
Rabr52 node_2 netRa52 -170927.31770803002
Lbr52 netRa52 netL52 -6.83276846198733e-11
Rbbr52 netL52 node_3 189068.00104529847
Cbr52 netL52 node_3 -2.116450636898347e-21

* Branch 53
Rabr53 node_2 netRa53 789749428.0114679
Lbr53 netRa53 netL53 2.609507240693683e-09
Rbbr53 netL53 node_3 -789777225.7331779
Cbr53 netL53 node_3 4.18376602188277e-27

* Branch 54
Rabr54 node_2 netRa54 894.4652695305502
Lbr54 netRa54 netL54 -1.8047745530839952e-11
Rbbr54 netL54 node_3 -409280.7026422536
Cbr54 netL54 node_3 -4.763473976967446e-20

* Branch 55
Rabr55 node_2 netRa55 -14299.840751223746
Lbr55 netRa55 netL55 -2.1253584367695297e-11
Rbbr55 netL55 node_3 118410.09946026295
Cbr55 netL55 node_3 -1.2584268282056396e-20

* Branch 56
Rabr56 node_2 netRa56 4939.503638424044
Lbr56 netRa56 netL56 -1.1901938157465348e-11
Rbbr56 netL56 node_3 -73001.16766923413
Cbr56 netL56 node_3 -3.288958708483007e-20

* Branch 57
Rabr57 node_2 netRa57 5106.10615636267
Lbr57 netRa57 netL57 -1.1182979021822098e-11
Rbbr57 netL57 node_3 -51834.22377481142
Cbr57 netL57 node_3 -4.213652962950615e-20

* Branch 58
Rabr58 node_2 netRa58 79986.75826658311
Lbr58 netRa58 netL58 -4.562228362733413e-11
Rbbr58 netL58 node_3 -118736.36857364871
Cbr58 netL58 node_3 -4.800499948890264e-21

* Branch 59
Rabr59 node_2 netRa59 4340826.770088787
Lbr59 netRa59 netL59 1.5575140859081907e-10
Rbbr59 netL59 node_3 -4360713.948251797
Cbr59 netL59 node_3 8.228402514596593e-24

* Branch 60
Rabr60 node_2 netRa60 -4996.357129809812
Lbr60 netRa60 netL60 -1.8221910944687306e-11
Rbbr60 netL60 node_3 160205.51871615602
Cbr60 netL60 node_3 -2.283208503742789e-20

* Branch 61
Rabr61 node_2 netRa61 -13591.055174399567
Lbr61 netRa61 netL61 -1.7502640731223386e-11
Rbbr61 netL61 node_3 40926.60887357014
Cbr61 netL61 node_3 -3.149247063074148e-20

* Branch 62
Rabr62 node_2 netRa62 -17032.425788352994
Lbr62 netRa62 netL62 -3.163902535618921e-11
Rbbr62 netL62 node_3 57121.323478697326
Cbr62 netL62 node_3 -3.2556255882946213e-20

* Branch 63
Rabr63 node_2 netRa63 -250639.03730932623
Lbr63 netRa63 netL63 -3.992955919770151e-11
Rbbr63 netL63 node_3 271951.4763815244
Cbr63 netL63 node_3 -5.858586802479468e-22

* Branch 64
Rabr64 node_2 netRa64 -48540.05004351919
Lbr64 netRa64 netL64 -2.8218392857184136e-11
Rbbr64 netL64 node_3 75916.58071997171
Cbr64 netL64 node_3 -7.659452609468265e-21

* Branch 65
Rabr65 node_2 netRa65 -26000.190801517052
Lbr65 netRa65 netL65 -4.0054663631265725e-11
Rbbr65 netL65 node_3 69924.7814159528
Cbr65 netL65 node_3 -2.2044767504231763e-20

* Branch 66
Rabr66 node_2 netRa66 -17622.980746901263
Lbr66 netRa66 netL66 -3.671055185829589e-11
Rbbr66 netL66 node_3 94941.71267007124
Cbr66 netL66 node_3 -2.19576130203959e-20

* Branch 67
Rabr67 node_2 netRa67 -8214.321671051775
Lbr67 netRa67 netL67 -5.770753765257097e-11
Rbbr67 netL67 node_3 403938.4309234362
Cbr67 netL67 node_3 -1.7425417585372202e-20

* Branch 68
Rabr68 node_2 netRa68 -31808.65147130347
Lbr68 netRa68 netL68 -3.849234522377028e-11
Rbbr68 netL68 node_3 67842.69758626226
Cbr68 netL68 node_3 -1.7842578129506225e-20

* Branch 69
Rabr69 node_2 netRa69 -22845.12386864232
Lbr69 netRa69 netL69 -3.194059344800859e-11
Rbbr69 netL69 node_3 69605.70687080798
Cbr69 netL69 node_3 -2.0092871103274134e-20

* Branch 70
Rabr70 node_2 netRa70 -38470.88184829327
Lbr70 netRa70 netL70 -4.0665826668145783e-11
Rbbr70 netL70 node_3 70379.51747287493
Cbr70 netL70 node_3 -1.50217622127146e-20

* Branch 71
Rabr71 node_2 netRa71 -41897.69781735246
Lbr71 netRa71 netL71 -4.020498412735531e-11
Rbbr71 netL71 node_3 72967.99633428175
Cbr71 netL71 node_3 -1.3152722118646544e-20

* Branch 72
Rabr72 node_2 netRa72 -38085.01764288183
Lbr72 netRa72 netL72 -3.350791676376993e-11
Rbbr72 netL72 node_3 62787.59304629972
Cbr72 netL72 node_3 -1.401427581648188e-20

* Branch 73
Rabr73 node_2 netRa73 -45780.834695093414
Lbr73 netRa73 netL73 -4.617730743143688e-11
Rbbr73 netL73 node_3 76171.64547626041
Cbr73 netL73 node_3 -1.3243428773872966e-20

* Branch 74
Rabr74 node_2 netRa74 34619.258688505084
Lbr74 netRa74 netL74 2.5574979889636294e-11
Rbbr74 netL74 node_3 -77618.06038969876
Cbr74 netL74 node_3 9.518505432435433e-21

* Branch 75
Rabr75 node_2 netRa75 -385054.0844082728
Lbr75 netRa75 netL75 -1.4596798042644584e-10
Rbbr75 netL75 node_3 414996.38454619196
Cbr75 netL75 node_3 -9.13496953762766e-22

* Branch 76
Rabr76 node_2 netRa76 -36544.77221366133
Lbr76 netRa76 netL76 -3.2875791527025035e-11
Rbbr76 netL76 node_3 96011.18081860957
Cbr76 netL76 node_3 -9.370317496550419e-21

* Branch 77
Rabr77 node_2 netRa77 -47040.69082427369
Lbr77 netRa77 netL77 -4.549504007686469e-11
Rbbr77 netL77 node_3 74490.0630740759
Cbr77 netL77 node_3 -1.2984267819845538e-20

* Branch 78
Rabr78 node_2 netRa78 -86965.32870585269
Lbr78 netRa78 netL78 -6.068424957682203e-11
Rbbr78 netL78 node_3 111028.97755358026
Cbr78 netL78 node_3 -6.284947259329092e-21

* Branch 79
Rabr79 node_2 netRa79 -65049.35416471811
Lbr79 netRa79 netL79 -5.2165462637710147e-11
Rbbr79 netL79 node_3 89971.27365793187
Cbr79 netL79 node_3 -8.913421131460019e-21

* Branch 80
Rabr80 node_2 netRa80 -40459.80632423402
Lbr80 netRa80 netL80 -3.0212365258071646e-11
Rbbr80 netL80 node_3 60097.32852288259
Cbr80 netL80 node_3 -1.242543931282813e-20

* Branch 81
Rabr81 node_2 netRa81 -22834.550445590314
Lbr81 netRa81 netL81 -4.0780776825540187e-11
Rbbr81 netL81 node_3 151337.99786149917
Cbr81 netL81 node_3 -1.1801220047515491e-20

* Branch 82
Rabr82 node_2 netRa82 -41845.13944475858
Lbr82 netRa82 netL82 -4.4296025841640936e-11
Rbbr82 netL82 node_3 92651.06710658489
Cbr82 netL82 node_3 -1.1425374101861594e-20

* Branch 83
Rabr83 node_2 netRa83 -19643.986106754764
Lbr83 netRa83 netL83 -2.580758703484438e-11
Rbbr83 netL83 node_3 57633.69881001635
Cbr83 netL83 node_3 -2.2795170219643634e-20

* Branch 84
Rabr84 node_2 netRa84 -56598.30823188331
Lbr84 netRa84 netL84 -4.106096681897565e-11
Rbbr84 netL84 node_3 70467.63959997997
Cbr84 netL84 node_3 -1.0295285019427175e-20

* Branch 85
Rabr85 node_2 netRa85 -12734.229307079342
Lbr85 netRa85 netL85 -1.653947133985363e-11
Rbbr85 netL85 node_3 57002.171060196204
Cbr85 netL85 node_3 -2.27863659638311e-20

* Branch 86
Rabr86 node_2 netRa86 55307.57119695776
Lbr86 netRa86 netL86 3.875142525882033e-11
Rbbr86 netL86 node_3 -66023.83825882286
Cbr86 netL86 node_3 1.0613003529852819e-20

* Branch 87
Rabr87 node_2 netRa87 -1592857.8455999827
Lbr87 netRa87 netL87 1.521145410714518e-10
Rbbr87 netL87 node_3 1600022.81076249
Cbr87 netL87 node_3 5.968419328725372e-23

* Branch 88
Rabr88 node_2 netRa88 2187926.696435874
Lbr88 netRa88 netL88 -2.234560523940588e-10
Rbbr88 netL88 node_3 -2222940.646768732
Cbr88 netL88 node_3 -4.594282842726236e-23

* Branch 89
Rabr89 node_2 netRa89 -214990.08552540472
Lbr89 netRa89 netL89 5.622202392089696e-11
Rbbr89 netL89 node_3 221502.95276097825
Cbr89 netL89 node_3 1.1805127394242641e-21

* Branch 90
Rabr90 node_2 netRa90 -16.155943251278707
Lbr90 netRa90 netL90 -1.1795060455448373e-11
Rbbr90 netL90 node_3 20843761.55576223
Cbr90 netL90 node_3 -4.680002465324979e-20

* Branch 91
Rabr91 node_2 netRa91 17529.186796999817
Lbr91 netRa91 netL91 -1.8921103447655854e-11
Rbbr91 netL91 node_3 -49754.281686176946
Cbr91 netL91 node_3 -2.1685597583480404e-20

* Branch 92
Rabr92 node_2 netRa92 882441.2675302126
Lbr92 netRa92 netL92 -1.3655336748557089e-10
Rbbr92 netL92 node_3 -908587.2880833531
Cbr92 netL92 node_3 -1.703002315372915e-22

* Branch 93
Rabr93 node_2 netRa93 46222.430982994454
Lbr93 netRa93 netL93 1.586046883436247e-11
Rbbr93 netL93 node_3 -61084.09661645912
Cbr93 netL93 node_3 5.618707156535763e-21

* Branch 94
Rabr94 node_2 netRa94 22896.276177212436
Lbr94 netRa94 netL94 -1.798291524304127e-11
Rbbr94 netL94 node_3 -62245.1240949826
Cbr94 netL94 node_3 -1.2610323169829842e-20

* Branch 95
Rabr95 node_2 netRa95 37746.24697779345
Lbr95 netRa95 netL95 -2.0940496856489004e-11
Rbbr95 netL95 node_3 -70813.64622094834
Cbr95 netL95 node_3 -7.830479492321985e-21

* Branch 96
Rabr96 node_2 netRa96 328995.4111073038
Lbr96 netRa96 netL96 -5.553229458289699e-11
Rbbr96 netL96 node_3 -340976.49662505765
Cbr96 netL96 node_3 -4.949543195635428e-22

* Branch 97
Rabr97 node_2 netRa97 95318.40046122011
Lbr97 netRa97 netL97 1.4707737036648582e-11
Rbbr97 netL97 node_3 -101390.22786007152
Cbr97 netL97 node_3 1.5221849942291078e-21

* Branch 98
Rabr98 node_2 netRa98 6185.428691851976
Lbr98 netRa98 netL98 -4.4998075965788135e-12
Rbbr98 netL98 node_3 -14736.818461002866
Cbr98 netL98 node_3 -4.927929729395369e-20

* Branch 99
Rabr99 node_2 netRa99 2111.2548514836144
Lbr99 netRa99 netL99 -1.91611413644393e-12
Rbbr99 netL99 node_3 -7137.973698113159
Cbr99 netL99 node_3 -1.2664637054702055e-19

.ends


* Y'24
.subckt yp24 node_2 node_4
* Branch 0
Rabr0 node_2 netRa0 1104.5277642889291
Lbr0 netRa0 netL0 -1.629826815822965e-12
Rbbr0 netL0 node_4 -7667.033167833989
Cbr0 netL0 node_4 -1.8050957077379552e-19

* Branch 1
Rabr1 node_2 netRa1 521.7965244644332
Lbr1 netRa1 netL1 -1.3311990346296252e-12
Rbbr1 netL1 node_4 -9438.822744587269
Cbr1 netL1 node_4 -2.4383754734229815e-19

* Branch 2
Rabr2 node_2 netRa2 -23.721373065074854
Lbr2 netRa2 netL2 -1.055015403513881e-12
Rbbr2 netL2 node_4 -183893.6049682569
Cbr2 netL2 node_4 -3.257615541041051e-19

* Branch 3
Rabr3 node_2 netRa3 267.9179335834657
Lbr3 netRa3 netL3 -5.588100935154647e-13
Rbbr3 netL3 node_4 -3448.1122906620294
Cbr3 netL3 node_4 -5.65070871908336e-19

* Branch 4
Rabr4 node_2 netRa4 -2084.361358614824
Lbr4 netRa4 netL4 8.261251386820104e-13
Rbbr4 netL4 node_4 3044.4614562493325
Cbr4 netL4 node_4 1.2870395059555957e-19

* Branch 5
Rabr5 node_2 netRa5 -11213.607820678815
Lbr5 netRa5 netL5 -2.917294738597008e-12
Rbbr5 netL5 node_4 13582.613474646816
Cbr5 netL5 node_4 -1.9296484514122535e-20

* Branch 6
Rabr6 node_2 netRa6 327506.5875042253
Lbr6 netRa6 netL6 -1.2023569613059137e-11
Rbbr6 netL6 node_4 -328622.68751649355
Cbr6 netL6 node_4 -1.1161795896380718e-22

* Branch 7
Rabr7 node_2 netRa7 40073.97455090473
Lbr7 netRa7 netL7 -5.767714118101429e-12
Rbbr7 netL7 node_4 -41773.917722358034
Cbr7 netL7 node_4 -3.433767232002642e-21

* Branch 8
Rabr8 node_2 netRa8 -1135.9842837486447
Lbr8 netRa8 netL8 1.5886385487082853e-12
Rbbr8 netL8 node_4 8114.060250222713
Cbr8 netL8 node_4 1.6696685655729502e-19

* Branch 9
Rabr9 node_2 netRa9 -495.2980829595056
Lbr9 netRa9 netL9 4.3464938280301713e-13
Rbbr9 netL9 node_4 1572.3920643511549
Cbr9 netL9 node_4 5.476836549434198e-19

* Branch 10
Rabr10 node_2 netRa10 323.52595621040666
Lbr10 netRa10 netL10 -4.4168392137437007e-13
Rbbr10 netL10 node_4 -1847.7296177610156
Cbr10 netL10 node_4 -7.189193606267242e-19

* Branch 11
Rabr11 node_2 netRa11 779.6728225199661
Lbr11 netRa11 netL11 -1.756532732407953e-12
Rbbr11 netL11 node_4 -9298.256741813462
Cbr11 netL11 node_4 -2.321250312773014e-19

* Branch 12
Rabr12 node_2 netRa12 71881.02932728313
Lbr12 netRa12 netL12 7.829324152816317e-12
Rbbr12 netL12 node_4 -73439.8285592954
Cbr12 netL12 node_4 1.4861237736329168e-21

* Branch 13
Rabr13 node_2 netRa13 2547.469269015962
Lbr13 netRa13 netL13 2.0787088126538296e-12
Rbbr13 netL13 node_4 -4783.735333543234
Cbr13 netL13 node_4 1.7318986006882913e-19

* Branch 14
Rabr14 node_2 netRa14 -2412.1784902041395
Lbr14 netRa14 netL14 1.7397686770608801e-12
Rbbr14 netL14 node_4 6434.124941412328
Cbr14 netL14 node_4 1.1062137401021542e-19

* Branch 15
Rabr15 node_2 netRa15 -968.0370918558773
Lbr15 netRa15 netL15 1.2353888344776294e-12
Rbbr15 netL15 node_4 5954.005094785014
Cbr15 netL15 node_4 2.0946950475190002e-19

* Branch 16
Rabr16 node_2 netRa16 3042.59004329508
Lbr16 netRa16 netL16 -7.14758561300739e-12
Rbbr16 netL16 node_4 -12259.853371589568
Cbr16 netL16 node_4 -1.8478830175419356e-19

* Branch 17
Rabr17 node_2 netRa17 -1300.8249375656947
Lbr17 netRa17 netL17 -3.4432000794526185e-12
Rbbr17 netL17 node_4 14303.215616575719
Cbr17 netL17 node_4 -1.9199468553793912e-19

* Branch 18
Rabr18 node_2 netRa18 -5075.635885418207
Lbr18 netRa18 netL18 2.3271999370569046e-12
Rbbr18 netL18 node_4 8749.041145814339
Cbr18 netL18 node_4 5.2107040266652004e-20

* Branch 19
Rabr19 node_2 netRa19 4579501.107832743
Lbr19 netRa19 netL19 1.1830599325365846e-10
Rbbr19 netL19 node_4 -4583621.929272937
Cbr19 netL19 node_4 5.63791776823057e-24

* Branch 20
Rabr20 node_2 netRa20 28146.924942634596
Lbr20 netRa20 netL20 5.844299325985056e-12
Rbbr20 netL20 node_4 -30488.899530432718
Cbr20 netL20 node_4 6.82725569152339e-21

* Branch 21
Rabr21 node_2 netRa21 67974.47488287541
Lbr21 netRa21 netL21 6.8491988640469765e-12
Rbbr21 netL21 node_4 -69489.7594877917
Cbr21 netL21 node_4 1.4517687118727786e-21

* Branch 22
Rabr22 node_2 netRa22 -6088178.210440046
Lbr22 netRa22 netL22 1.2767315306750255e-10
Rbbr22 netL22 node_4 6093169.819060501
Cbr22 netL22 node_4 3.4408286666902724e-24

* Branch 23
Rabr23 node_2 netRa23 -45636.06649091213
Lbr23 netRa23 netL23 -9.24443975672956e-12
Rbbr23 netL23 node_4 49334.60487340814
Cbr23 netL23 node_4 -4.1156884680216345e-21

* Branch 24
Rabr24 node_2 netRa24 5967.384263149607
Lbr24 netRa24 netL24 -4.746980870342151e-12
Rbbr24 netL24 node_4 -8768.681807073648
Cbr24 netL24 node_4 -8.989502397846099e-20

* Branch 25
Rabr25 node_2 netRa25 197.32554477674032
Lbr25 netRa25 netL25 8.356261424370435e-13
Rbbr25 netL25 node_4 -9187.3459353553
Cbr25 netL25 node_4 4.84188098618894e-19

* Branch 26
Rabr26 node_2 netRa26 520571.6912232087
Lbr26 netRa26 netL26 -2.73545508897097e-11
Rbbr26 netL26 node_4 -522214.87313035334
Cbr26 netL26 node_4 -1.0056520166399197e-22

* Branch 27
Rabr27 node_2 netRa27 1042652.7382155594
Lbr27 netRa27 netL27 -4.044257538402872e-11
Rbbr27 netL27 node_4 -1044030.4894854167
Cbr27 netL27 node_4 -3.713644729977209e-23

* Branch 28
Rabr28 node_2 netRa28 11057.701578641609
Lbr28 netRa28 netL28 -3.794749925469897e-12
Rbbr28 netL28 node_4 -13107.248247541618
Cbr28 netL28 node_4 -2.6085868724346546e-20

* Branch 29
Rabr29 node_2 netRa29 -105.66095838381418
Lbr29 netRa29 netL29 1.08693607599896e-12
Rbbr29 netL29 node_4 21860.600765758292
Cbr29 netL29 node_4 4.2366658111119706e-19

* Branch 30
Rabr30 node_2 netRa30 5719.732655730846
Lbr30 netRa30 netL30 -4.389943057114426e-12
Rbbr30 netL30 node_4 -9065.222649544266
Cbr30 netL30 node_4 -8.398748699087575e-20

* Branch 31
Rabr31 node_2 netRa31 104703.50534268202
Lbr31 netRa31 netL31 -9.631394945436043e-12
Rbbr31 netL31 node_4 -106877.05594973128
Cbr31 netL31 node_4 -8.598621017079845e-22

* Branch 32
Rabr32 node_2 netRa32 8179.196796660482
Lbr32 netRa32 netL32 -4.576404636211816e-12
Rbbr32 netL32 node_4 -10834.847034690603
Cbr32 netL32 node_4 -5.1346315072375476e-20

* Branch 33
Rabr33 node_2 netRa33 -2257.076638792264
Lbr33 netRa33 netL33 -1.4730134834388193e-12
Rbbr33 netL33 node_4 5330.48650053421
Cbr33 netL33 node_4 -1.2325172473040585e-19

* Branch 34
Rabr34 node_2 netRa34 2675.9547779815757
Lbr34 netRa34 netL34 6.488784891999935e-13
Rbbr34 netL34 node_4 -3119.0962226615993
Cbr34 netL34 node_4 7.792051317157918e-20

* Branch 35
Rabr35 node_2 netRa35 -21497.504211815165
Lbr35 netRa35 netL35 -3.839594637099945e-12
Rbbr35 netL35 node_4 23335.19468511694
Cbr35 netL35 node_4 -7.666635151768703e-21

* Branch 36
Rabr36 node_2 netRa36 10067.970728529426
Lbr36 netRa36 netL36 -5.139404462980553e-12
Rbbr36 netL36 node_4 -12202.717463264189
Cbr36 netL36 node_4 -4.164114208155467e-20

* Branch 37
Rabr37 node_2 netRa37 -3072.1269761082826
Lbr37 netRa37 netL37 -7.31608677322982e-12
Rbbr37 netL37 node_4 19471.338445141686
Cbr37 netL37 node_4 -1.248332920103719e-19

* Branch 38
Rabr38 node_2 netRa38 3121.649122838576
Lbr38 netRa38 netL38 -5.736866735093443e-12
Rbbr38 netL38 node_4 -9308.655847297587
Cbr38 netL38 node_4 -1.9459327161209751e-19

* Branch 39
Rabr39 node_2 netRa39 1075.4863777343523
Lbr39 netRa39 netL39 -2.5984806643476594e-12
Rbbr39 netL39 node_4 -11699.6119363502
Cbr39 netL39 node_4 -2.0282644568888846e-19

* Branch 40
Rabr40 node_2 netRa40 -1225.6415318200488
Lbr40 netRa40 netL40 -2.626465993301636e-12
Rbbr40 netL40 node_4 10575.743049432334
Cbr40 netL40 node_4 -2.0580012931877383e-19

* Branch 41
Rabr41 node_2 netRa41 42405.36101867972
Lbr41 netRa41 netL41 -4.857980833808372e-12
Rbbr41 netL41 node_4 -43688.07785374701
Cbr41 netL41 node_4 -2.6201456303523194e-21

* Branch 42
Rabr42 node_2 netRa42 6850.799186957717
Lbr42 netRa42 netL42 -3.15173071064155e-12
Rbbr42 netL42 node_4 -9103.287777408384
Cbr42 netL42 node_4 -5.0385147217540475e-20

* Branch 43
Rabr43 node_2 netRa43 2105.239135003988
Lbr43 netRa43 netL43 -2.7391338879472495e-12
Rbbr43 netL43 node_4 -7285.402522278588
Cbr43 netL43 node_4 -1.7708411854559473e-19

* Branch 44
Rabr44 node_2 netRa44 1904.6488198195973
Lbr44 netRa44 netL44 2.6767912834408376e-12
Rbbr44 netL44 node_4 -7394.326605676783
Cbr44 netL44 node_4 1.9175916921171245e-19

* Branch 45
Rabr45 node_2 netRa45 2671.3259095530057
Lbr45 netRa45 netL45 -1.154665495955323e-12
Rbbr45 netL45 node_4 -4095.4523669365162
Cbr45 netL45 node_4 -1.0527437200026737e-19

* Branch 46
Rabr46 node_2 netRa46 -1138339.1615642037
Lbr46 netRa46 netL46 -9.696937711414963e-11
Rbbr46 netL46 node_4 1146132.8692960571
Cbr46 netL46 node_4 -7.436085851730661e-23

* Branch 47
Rabr47 node_2 netRa47 -7529.728721433097
Lbr47 netRa47 netL47 7.2248387806241054e-12
Rbbr47 netL47 node_4 17229.7012970816
Cbr47 netL47 node_4 5.540794358180641e-20

* Branch 48
Rabr48 node_2 netRa48 -24279.972113760436
Lbr48 netRa48 netL48 -4.209590824819052e-12
Rbbr48 netL48 node_4 26278.711689659114
Cbr48 netL48 node_4 -6.603359152495414e-21

* Branch 49
Rabr49 node_2 netRa49 788.9948464244441
Lbr49 netRa49 netL49 2.1684716522308323e-12
Rbbr49 netL49 node_4 -11143.856098381166
Cbr49 netL49 node_4 2.499457906717099e-19

* Branch 50
Rabr50 node_2 netRa50 -777668.7028278137
Lbr50 netRa50 netL50 -5.500165360491504e-11
Rbbr50 netL50 node_4 783481.9461157843
Cbr50 netL50 node_4 -9.030084649435338e-23

* Branch 51
Rabr51 node_2 netRa51 40625.68879318833
Lbr51 netRa51 netL51 1.0555300832221126e-11
Rbbr51 netL51 node_4 -49637.55584204604
Cbr51 netL51 node_4 5.2404195639343005e-21

* Branch 52
Rabr52 node_2 netRa52 -17761.346222957105
Lbr52 netRa52 netL52 1.1284591501514269e-11
Rbbr52 netL52 node_4 21494.72094050787
Cbr52 netL52 node_4 2.948506533140699e-20

* Branch 53
Rabr53 node_2 netRa53 -29416.39202704677
Lbr53 netRa53 netL53 8.25634526950571e-12
Rbbr53 netL53 node_4 34932.750542885515
Cbr53 netL53 node_4 8.026254107090937e-21

* Branch 54
Rabr54 node_2 netRa54 -3378.1435712929347
Lbr54 netRa54 netL54 4.659148403592135e-12
Rbbr54 netL54 node_4 11079.742915033905
Cbr54 netL54 node_4 1.238450300619579e-19

* Branch 55
Rabr55 node_2 netRa55 -11863.112109138296
Lbr55 netRa55 netL55 7.356395476687119e-12
Rbbr55 netL55 node_4 21485.756836623827
Cbr55 netL55 node_4 2.8801719753218036e-20

* Branch 56
Rabr56 node_2 netRa56 -19191.62663922817
Lbr56 netRa56 netL56 6.6560844537013725e-12
Rbbr56 netL56 node_4 23612.82836040956
Cbr56 netL56 node_4 1.4671748508834874e-20

* Branch 57
Rabr57 node_2 netRa57 252.26868051457066
Lbr57 netRa57 netL57 -3.2602024418418444e-12
Rbbr57 netL57 node_4 -18201.987790700085
Cbr57 netL57 node_4 -6.836785256212962e-19

* Branch 58
Rabr58 node_2 netRa58 53399.50601315262
Lbr58 netRa58 netL58 1.0621334052499728e-11
Rbbr58 netL58 node_4 -60469.02602234573
Cbr58 netL58 node_4 3.29128172260615e-21

* Branch 59
Rabr59 node_2 netRa59 5644.877344393285
Lbr59 netRa59 netL59 -5.363517545472249e-12
Rbbr59 netL59 node_4 -9025.136384192423
Cbr59 netL59 node_4 -1.05008719825373e-19

* Branch 60
Rabr60 node_2 netRa60 -2467039.9096712973
Lbr60 netRa60 netL60 1.2434276196047655e-10
Rbbr60 netL60 node_4 2474784.505080657
Cbr60 netL60 node_4 2.03633640287192e-23

* Branch 61
Rabr61 node_2 netRa61 -14132644.598897919
Lbr61 netRa61 netL61 -3.6407823546133666e-10
Rbbr61 netL61 node_4 14143553.739949873
Cbr61 netL61 node_4 -1.8215537954454152e-24

* Branch 62
Rabr62 node_2 netRa62 218901.96825362064
Lbr62 netRa62 netL62 7.651019420358573e-11
Rbbr62 netL62 node_4 -232049.1104695729
Cbr62 netL62 node_4 1.5073797060180197e-21

* Branch 63
Rabr63 node_2 netRa63 -92608.76025806012
Lbr63 netRa63 netL63 -2.3975690966370873e-11
Rbbr63 netL63 node_4 107083.86085402376
Cbr63 netL63 node_4 -2.4190056014567566e-21

* Branch 64
Rabr64 node_2 netRa64 -55552.88059714492
Lbr64 netRa64 netL64 -6.127547252569854e-12
Rbbr64 netL64 node_4 57440.11229978085
Cbr64 netL64 node_4 -1.9206867742621223e-21

* Branch 65
Rabr65 node_2 netRa65 -17856.057222547082
Lbr65 netRa65 netL65 -5.123403426170212e-12
Rbbr65 netL65 node_4 21706.15380198745
Cbr65 netL65 node_4 -1.3225258176813326e-20

* Branch 66
Rabr66 node_2 netRa66 99.08798836621317
Lbr66 netRa66 netL66 1.2753852683818727e-11
Rbbr66 netL66 node_4 -1345892.3084495633
Cbr66 netL66 node_4 1.1503291818700914e-19

* Branch 67
Rabr67 node_2 netRa67 -482227.08162364434
Lbr67 netRa67 netL67 5.885149010089688e-11
Rbbr67 netL67 node_4 507761.2956389207
Cbr67 netL67 node_4 2.4031516351995045e-22

* Branch 68
Rabr68 node_2 netRa68 -50609.78171889758
Lbr68 netRa68 netL68 3.636886476221461e-11
Rbbr68 netL68 node_4 76084.59602913701
Cbr68 netL68 node_4 9.438056710455267e-21

* Branch 69
Rabr69 node_2 netRa69 1786.610970205543
Lbr69 netRa69 netL69 1.1526677197114363e-11
Rbbr69 netL69 node_4 -85654.62367462824
Cbr69 netL69 node_4 7.578032056134915e-20

* Branch 70
Rabr70 node_2 netRa70 3687.110564847488
Lbr70 netRa70 netL70 1.7091010553290472e-11
Rbbr70 netL70 node_4 -60282.11739030245
Cbr70 netL70 node_4 7.719365253635587e-20

* Branch 71
Rabr71 node_2 netRa71 -29008.26733099502
Lbr71 netRa71 netL71 -9.735232383317873e-12
Rbbr71 netL71 node_4 36452.02086840308
Cbr71 netL71 node_4 -9.208739923612236e-21

* Branch 72
Rabr72 node_2 netRa72 -2594.516103021
Lbr72 netRa72 netL72 1.6540300534878915e-11
Rbbr72 netL72 node_4 108717.45815522996
Cbr72 netL72 node_4 5.840639270680038e-20

* Branch 73
Rabr73 node_2 netRa73 5764.108984985478
Lbr73 netRa73 netL73 1.7995177343146455e-11
Rbbr73 netL73 node_4 -49288.10200159784
Cbr73 netL73 node_4 6.344760311367849e-20

* Branch 74
Rabr74 node_2 netRa74 5178.521388019915
Lbr74 netRa74 netL74 9.281702288887625e-12
Rbbr74 netL74 node_4 -19672.610950153074
Cbr74 netL74 node_4 9.11883136406685e-20

* Branch 75
Rabr75 node_2 netRa75 592.1700425760565
Lbr75 netRa75 netL75 2.428246851835846e-11
Rbbr75 netL75 node_4 -1100085.1298617146
Cbr75 netL75 node_4 3.7979461697844874e-20

* Branch 76
Rabr76 node_2 netRa76 684.1115044892771
Lbr76 netRa76 netL76 1.3206004762674412e-11
Rbbr76 netL76 node_4 -269826.77583583636
Cbr76 netL76 node_4 7.215750069730316e-20

* Branch 77
Rabr77 node_2 netRa77 10323.31701843208
Lbr77 netRa77 netL77 1.662437892809869e-11
Rbbr77 netL77 node_4 -31895.86933832063
Cbr77 netL77 node_4 5.0522251785214887e-20

* Branch 78
Rabr78 node_2 netRa78 7967.294406459714
Lbr78 netRa78 netL78 1.576021202834068e-11
Rbbr78 netL78 node_4 -34104.73699560978
Cbr78 netL78 node_4 5.804225230292149e-20

* Branch 79
Rabr79 node_2 netRa79 11335.658743119606
Lbr79 netRa79 netL79 1.8273632310369822e-11
Rbbr79 netL79 node_4 -33210.55414694547
Cbr79 netL79 node_4 4.856576130221146e-20

* Branch 80
Rabr80 node_2 netRa80 21153.162530808404
Lbr80 netRa80 netL80 2.6239897547079935e-11
Rbbr80 netL80 node_4 -42394.37558550453
Cbr80 netL80 node_4 2.9268404739236534e-20

* Branch 81
Rabr81 node_2 netRa81 474679.909428157
Lbr81 netRa81 netL81 1.6570496630032914e-10
Rbbr81 netL81 node_4 -506004.74290927936
Cbr81 netL81 node_4 6.899259446845179e-22

* Branch 82
Rabr82 node_2 netRa82 20198.753926523168
Lbr82 netRa82 netL82 2.6920035108205276e-11
Rbbr82 netL82 node_4 -42582.543001570964
Cbr82 netL82 node_4 3.130328015674229e-20

* Branch 83
Rabr83 node_2 netRa83 31834.778542532473
Lbr83 netRa83 netL83 2.945412053513611e-11
Rbbr83 netL83 node_4 -48069.29837831483
Cbr83 netL83 node_4 1.924874552256466e-20

* Branch 84
Rabr84 node_2 netRa84 86333.10250884457
Lbr84 netRa84 netL84 5.0692609308903325e-11
Rbbr84 netL84 node_4 -103248.10749993943
Cbr84 netL84 node_4 5.687218790687877e-21

* Branch 85
Rabr85 node_2 netRa85 353134.324009201
Lbr85 netRa85 netL85 -3.048224539230964e-11
Rbbr85 netL85 node_4 -356349.6422115214
Cbr85 netL85 node_4 -2.422314231463267e-22

* Branch 86
Rabr86 node_2 netRa86 32842.549234328784
Lbr86 netRa86 netL86 2.979449914945429e-11
Rbbr86 netL86 node_4 -45428.69094005409
Cbr86 netL86 node_4 1.9969924579701243e-20

* Branch 87
Rabr87 node_2 netRa87 46095.14200892484
Lbr87 netRa87 netL87 3.065047667621327e-11
Rbbr87 netL87 node_4 -80126.80331329527
Cbr87 netL87 node_4 8.299046298392285e-21

* Branch 88
Rabr88 node_2 netRa88 873.1214446295014
Lbr88 netRa88 netL88 4.297566083006676e-11
Rbbr88 netL88 node_4 -4385999.935051747
Cbr88 netL88 node_4 1.1280634798237286e-20

* Branch 89
Rabr89 node_2 netRa89 221.24364757076756
Lbr89 netRa89 netL89 -8.001652405491006e-12
Rbbr89 netL89 node_4 -143570.90656270206
Cbr89 netL89 node_4 -2.503784422237722e-19

* Branch 90
Rabr90 node_2 netRa90 23492.79261844038
Lbr90 netRa90 netL90 2.548290471386604e-11
Rbbr90 netL90 node_4 -79086.37205162049
Cbr90 netL90 node_4 1.3718150750388703e-20

* Branch 91
Rabr91 node_2 netRa91 -16346.659174226621
Lbr91 netRa91 netL91 -1.7850150004778013e-11
Rbbr91 netL91 node_4 24040.798913579434
Cbr91 netL91 node_4 -4.543525339304223e-20

* Branch 92
Rabr92 node_2 netRa92 -112577.84366003214
Lbr92 netRa92 netL92 6.279616479848512e-11
Rbbr92 netL92 node_4 166313.03350338928
Cbr92 netL92 node_4 3.3534115870696332e-21

* Branch 93
Rabr93 node_2 netRa93 -1706.5655476011445
Lbr93 netRa93 netL93 2.6340576437451228e-12
Rbbr93 netL93 node_4 3518.9060010670432
Cbr93 netL93 node_4 4.384056464130499e-19

* Branch 94
Rabr94 node_2 netRa94 -24969.311282965566
Lbr94 netRa94 netL94 3.044811455765104e-11
Rbbr94 netL94 node_4 90455.89170050429
Cbr94 netL94 node_4 1.3475174425778396e-20

* Branch 95
Rabr95 node_2 netRa95 -2304.973688837727
Lbr95 netRa95 netL95 6.131141321566715e-12
Rbbr95 netL95 node_4 28014.744667216153
Cbr95 netL95 node_4 9.48539893085668e-20

* Branch 96
Rabr96 node_2 netRa96 -5553.143911936562
Lbr96 netRa96 netL96 -1.54862157555318e-11
Rbbr96 netL96 node_4 144974.37631215723
Cbr96 netL96 node_4 -1.926191373282477e-20

* Branch 97
Rabr97 node_2 netRa97 -10326.674022913276
Lbr97 netRa97 netL97 1.2073029078350663e-11
Rbbr97 netL97 node_4 28355.936955598867
Cbr97 netL97 node_4 4.1203629736956716e-20

* Branch 98
Rabr98 node_2 netRa98 -2586.2902741975267
Lbr98 netRa98 netL98 7.345540798185709e-12
Rbbr98 netL98 node_4 40316.442085329414
Cbr98 netL98 node_4 7.033023785274596e-20

* Branch 99
Rabr99 node_2 netRa99 -631.9330484912855
Lbr99 netRa99 netL99 -8.476077545766396e-13
Rbbr99 netL99 node_4 4098.26778225125
Cbr99 netL99 node_4 -3.432637140711891e-19

.ends


* Y'33
.subckt yp33 node_3 0
* Branch 0
Rabr0 node_3 netRa0 -8528794.802240271
Lbr0 netRa0 netL0 1.6433384475778716e-09
Rbbr0 netL0 0 9129768.203938976
Cbr0 netL0 0 2.1010228861773916e-23

* Branch 1
Rabr1 node_3 netRa1 -379602.3882159107
Lbr1 netRa1 netL1 1.1904515923450025e-10
Rbbr1 netL1 0 509080.5472669613
Cbr1 netL1 0 6.117892584778741e-22

* Branch 2
Rabr2 node_3 netRa2 2289377.99347533
Lbr2 netRa2 netL2 2.31143429934768e-09
Rbbr2 netL2 0 -7012012.659154626
Cbr2 netL2 0 1.4723284507250657e-22

* Branch 3
Rabr3 node_3 netRa3 57065.87056367981
Lbr3 netRa3 netL3 2.2123788550896239e-10
Rbbr3 netL3 0 -2563017.4257995132
Cbr3 netL3 0 1.641462542966423e-21

* Branch 4
Rabr4 node_3 netRa4 -1188725.5289051554
Lbr4 netRa4 netL4 1.9994314320807027e-10
Rbbr4 netL4 0 1305912.928642172
Cbr4 netL4 0 1.2840505273268335e-22

* Branch 5
Rabr5 node_3 netRa5 -5083131.122464335
Lbr5 netRa5 netL5 -5.42240519085027e-10
Rbbr5 netL5 0 5286214.171556748
Cbr5 netL5 0 -2.0211379524345808e-23

* Branch 6
Rabr6 node_3 netRa6 140150.5711654079
Lbr6 netRa6 netL6 6.123587116991671e-10
Rbbr6 netL6 0 -6630867.409719073
Cbr6 netL6 0 7.037193850726802e-22

* Branch 7
Rabr7 node_3 netRa7 -168037.70213668127
Lbr7 netRa7 netL7 2.903669316274984e-10
Rbbr7 netL7 0 1364732.434675781
Cbr7 netL7 0 1.2362058139374622e-21

* Branch 8
Rabr8 node_3 netRa8 -95943.92868929135
Lbr8 netRa8 netL8 4.745118358891781e-10
Rbbr8 netL8 0 4082544.9018526147
Cbr8 netL8 0 1.1352455990202747e-21

* Branch 9
Rabr9 node_3 netRa9 86659.10955901403
Lbr9 netRa9 netL9 8.09477785546462e-10
Rbbr9 netL9 0 -9886407.663293019
Cbr9 netL9 0 1.0692962083799506e-21

* Branch 10
Rabr10 node_3 netRa10 91113.89737606511
Lbr10 netRa10 netL10 8.06073683956384e-10
Rbbr10 netL10 0 -8609070.73842137
Cbr10 netL10 0 1.140869416687094e-21

* Branch 11
Rabr11 node_3 netRa11 19053.947733972283
Lbr11 netRa11 netL11 6.443074192133339e-10
Rbbr11 netL11 0 -57125713.22692625
Cbr11 netL11 0 9.533008972135322e-22

* Branch 12
Rabr12 node_3 netRa12 82209.86100297146
Lbr12 netRa12 netL12 7.877274036676185e-10
Rbbr12 netL12 0 -10491483.957806634
Cbr12 netL12 0 1.0199590374031493e-21

* Branch 13
Rabr13 node_3 netRa13 196162.74226730526
Lbr13 netRa13 netL13 1.874609893681125e-09
Rbbr13 netL13 0 -13999779.432051387
Cbr13 netL13 0 7.615467206449565e-22

* Branch 14
Rabr14 node_3 netRa14 816087.8518891562
Lbr14 netRa14 netL14 3.7514087290059165e-10
Rbbr14 netL14 0 -1355778.4717997606
Cbr14 netL14 0 3.4072409290862776e-22

* Branch 15
Rabr15 node_3 netRa15 185851.16056121685
Lbr15 netRa15 netL15 6.411914169562937e-10
Rbbr15 netL15 0 -5235678.37820951
Cbr15 netL15 0 6.817090006701363e-22

* Branch 16
Rabr16 node_3 netRa16 52213.162425982984
Lbr16 netRa16 netL16 6.832752327093322e-10
Rbbr16 netL16 0 -15555146.452868193
Cbr16 netL16 0 9.59060276908662e-22

* Branch 17
Rabr17 node_3 netRa17 81292.03596495911
Lbr17 netRa17 netL17 7.681975553372646e-10
Rbbr17 netL17 0 -10657827.041100642
Cbr17 netL17 0 9.724959204565013e-22

* Branch 18
Rabr18 node_3 netRa18 435942.5019714224
Lbr18 netRa18 netL18 8.196839130959836e-10
Rbbr18 netL18 0 -3695019.929522534
Cbr18 netL18 0 5.179018356287627e-22

* Branch 19
Rabr19 node_3 netRa19 58036.29461763318
Lbr19 netRa19 netL19 7.185197086852087e-10
Rbbr19 netL19 0 -14483251.595536573
Cbr19 netL19 0 9.6483228429444e-22

* Branch 20
Rabr20 node_3 netRa20 220199.62462146307
Lbr20 netRa20 netL20 7.407603363208375e-10
Rbbr20 netL20 0 -2528684.969926263
Cbr20 netL20 0 1.3719296174152006e-21

* Branch 21
Rabr21 node_3 netRa21 15634125.785411298
Lbr21 netRa21 netL21 -2.0839276000206058e-08
Rbbr21 netL21 0 -36202662.449828625
Cbr21 netL21 0 -3.647529455505376e-23

* Branch 22
Rabr22 node_3 netRa22 -1241.976359696673
Lbr22 netRa22 netL22 2.017230153605395e-10
Rbbr22 netL22 0 9151522.416481998
Cbr22 netL22 0 8.289353380551994e-21

* Branch 23
Rabr23 node_3 netRa23 220830.87426585783
Lbr23 netRa23 netL23 1.6263171737948625e-09
Rbbr23 netL23 0 -6303393.133059297
Cbr23 netL23 0 1.2298924277656533e-21

* Branch 24
Rabr24 node_3 netRa24 286183.7480787786
Lbr24 netRa24 netL24 -1.4109105309531285e-10
Rbbr24 netL24 0 -459009.66656128236
Cbr24 netL24 0 -1.070638902746007e-21

* Branch 25
Rabr25 node_3 netRa25 862454.2661789197
Lbr25 netRa25 netL25 1.8423402449292606e-09
Rbbr25 netL25 0 -3050839.3779228358
Cbr25 netL25 0 7.096484792518326e-22

* Branch 26
Rabr26 node_3 netRa26 93578.48012369146
Lbr26 netRa26 netL26 7.855816974799042e-10
Rbbr26 netL26 0 -6897807.717578116
Cbr26 netL26 0 1.283226327462312e-21

* Branch 27
Rabr27 node_3 netRa27 232038.30772201004
Lbr27 netRa27 netL27 4.97718046374007e-10
Rbbr27 netL27 0 -1135472.1518907936
Cbr27 netL27 0 1.9106185218138738e-21

* Branch 28
Rabr28 node_3 netRa28 -11803.851597661112
Lbr28 netRa28 netL28 -6.940381144322759e-11
Rbbr28 netL28 0 1217331.2179760365
Cbr28 netL28 0 -4.972228429052333e-21

* Branch 29
Rabr29 node_3 netRa29 2599064.872464191
Lbr29 netRa29 netL29 6.692832608080145e-10
Rbbr29 netL29 0 -2738492.2143846564
Cbr29 netL29 0 9.414772769751626e-23

* Branch 30
Rabr30 node_3 netRa30 -24045.56989714333
Lbr30 netRa30 netL30 8.482113310307006e-11
Rbbr30 netL30 0 851486.8136398299
Cbr30 netL30 0 4.0831691177052495e-21

* Branch 31
Rabr31 node_3 netRa31 126920.45786012732
Lbr31 netRa31 netL31 -1.318700987787639e-10
Rbbr31 netL31 0 -483818.6626383846
Cbr31 netL31 0 -2.1392337748537048e-21

* Branch 32
Rabr32 node_3 netRa32 -2640.0665092781705
Lbr32 netRa32 netL32 1.0254474245328449e-10
Rbbr32 netL32 0 9761574.04950693
Cbr32 netL32 0 3.501556894298904e-21

* Branch 33
Rabr33 node_3 netRa33 5015994.609475601
Lbr33 netRa33 netL33 -1.3081997120704761e-09
Rbbr33 netL33 0 -6045107.453625684
Cbr33 netL33 0 -4.310712193249571e-23

* Branch 34
Rabr34 node_3 netRa34 776957.351270619
Lbr34 netRa34 netL34 4.5606903691412566e-10
Rbbr34 netL34 0 -984790.4167989228
Cbr34 netL34 0 5.970873168321006e-22

* Branch 35
Rabr35 node_3 netRa35 -20402.05060981284
Lbr35 netRa35 netL35 5.351817706779165e-10
Rbbr35 netL35 0 22952018.195186578
Cbr35 netL35 0 1.0670902615726081e-21

* Branch 36
Rabr36 node_3 netRa36 -11284272.48823005
Lbr36 netRa36 netL36 1.6939538693809246e-09
Rbbr36 netL36 0 11442204.885456035
Cbr36 netL36 0 1.3114361174375893e-23

* Branch 37
Rabr37 node_3 netRa37 1765749.3000517942
Lbr37 netRa37 netL37 -3.3890542289453734e-10
Rbbr37 netL37 0 -1967277.0853506173
Cbr37 netL37 0 -9.751931376481577e-23

* Branch 38
Rabr38 node_3 netRa38 -1599069.4861904955
Lbr38 netRa38 netL38 -4.590794905319446e-10
Rbbr38 netL38 0 1924301.1634604305
Cbr38 netL38 0 -1.492885536992644e-22

* Branch 39
Rabr39 node_3 netRa39 88589.97260517816
Lbr39 netRa39 netL39 -2.9140533125727163e-10
Rbbr39 netL39 0 -685206.5882684382
Cbr39 netL39 0 -4.769867067010782e-21

* Branch 40
Rabr40 node_3 netRa40 114339.25785545295
Lbr40 netRa40 netL40 1.4609729022953685e-10
Rbbr40 netL40 0 -682886.9310646922
Cbr40 netL40 0 1.8745142873431676e-21

* Branch 41
Rabr41 node_3 netRa41 779866.4105499221
Lbr41 netRa41 netL41 -1.3893256681798417e-10
Rbbr41 netL41 0 -864795.0213697668
Cbr41 netL41 0 -2.0595150031003832e-22

* Branch 42
Rabr42 node_3 netRa42 127009.90022430681
Lbr42 netRa42 netL42 3.2099153576648955e-10
Rbbr42 netL42 0 -809777.0150901757
Cbr42 netL42 0 3.13095017409624e-21

* Branch 43
Rabr43 node_3 netRa43 64134.658938315966
Lbr43 netRa43 netL43 1.86072759414841e-10
Rbbr43 netL43 0 -1845227.8951732875
Cbr43 netL43 0 1.5780082547019436e-21

* Branch 44
Rabr44 node_3 netRa44 114201.78649204
Lbr44 netRa44 netL44 -4.445224085381987e-10
Rbbr44 netL44 0 -1237651.5618808568
Cbr44 netL44 0 -3.13203294828478e-21

* Branch 45
Rabr45 node_3 netRa45 145550.20682227024
Lbr45 netRa45 netL45 -1.8394395427255716e-10
Rbbr45 netL45 0 -821433.0700921165
Cbr45 netL45 0 -1.537217735635028e-21

* Branch 46
Rabr46 node_3 netRa46 2745.397069668743
Lbr46 netRa46 netL46 3.4560950076867977e-10
Rbbr46 netL46 0 -41297307.408912174
Cbr46 netL46 0 3.1907245989004652e-21

* Branch 47
Rabr47 node_3 netRa47 -89400.24385196215
Lbr47 netRa47 netL47 7.531875136598087e-10
Rbbr47 netL47 0 5606252.078247678
Cbr47 netL47 0 1.498653084483082e-21

* Branch 48
Rabr48 node_3 netRa48 426363.47350524244
Lbr48 netRa48 netL48 -1.074363413033565e-09
Rbbr48 netL48 0 -2270188.8449741416
Cbr48 netL48 0 -1.1091181995069236e-21

* Branch 49
Rabr49 node_3 netRa49 2907890.5095284646
Lbr49 netRa49 netL49 -6.342158668673535e-10
Rbbr49 netL49 0 -3230257.60190619
Cbr49 netL49 0 -6.751407560010529e-23

* Branch 50
Rabr50 node_3 netRa50 -417048.38627957576
Lbr50 netRa50 netL50 7.907827276249735e-10
Rbbr50 netL50 0 2521807.341183117
Cbr50 netL50 0 7.515593512872185e-22

* Branch 51
Rabr51 node_3 netRa51 1243149.1929299908
Lbr51 netRa51 netL51 2.1203960180523394e-09
Rbbr51 netL51 0 -3300275.8383047106
Cbr51 netL51 0 5.170213406947184e-22

* Branch 52
Rabr52 node_3 netRa52 5314898.896929072
Lbr52 netRa52 netL52 3.4450803480931232e-09
Rbbr52 netL52 0 -6525017.421035834
Cbr52 netL52 0 9.934961874607078e-23

* Branch 53
Rabr53 node_3 netRa53 2576002.1314337007
Lbr53 netRa53 netL53 -4.703671976843905e-10
Rbbr53 netL53 0 -2853018.478503439
Cbr53 netL53 0 -6.39992953059597e-23

* Branch 54
Rabr54 node_3 netRa54 41970504.05304379
Lbr54 netRa54 netL54 8.347934984679535e-09
Rbbr54 netL54 0 -42784701.80451452
Cbr54 netL54 0 4.6489873248249044e-24

* Branch 55
Rabr55 node_3 netRa55 4366564.033171941
Lbr55 netRa55 netL55 3.0648303314832218e-09
Rbbr55 netL55 0 -5476196.987235654
Cbr55 netL55 0 1.2818264633496227e-22

* Branch 56
Rabr56 node_3 netRa56 45845944.9005491
Lbr56 netRa56 netL56 -1.1369517504963931e-08
Rbbr56 netL56 0 -47853349.86904291
Cbr56 netL56 0 -5.182209646050531e-24

* Branch 57
Rabr57 node_3 netRa57 -365766.7213756204
Lbr57 netRa57 netL57 8.771228618691761e-10
Rbbr57 netL57 0 4280287.193616887
Cbr57 netL57 0 5.601036897899676e-22

* Branch 58
Rabr58 node_3 netRa58 403899.30177527555
Lbr58 netRa58 netL58 -1.5359308537200098e-09
Rbbr58 netL58 0 -4738377.695334366
Cbr58 netL58 0 -8.022430391892085e-22

* Branch 59
Rabr59 node_3 netRa59 -4653249.63306671
Lbr59 netRa59 netL59 2.101854878522877e-09
Rbbr59 netL59 0 6110238.591718782
Cbr59 netL59 0 7.39212260731016e-23

* Branch 60
Rabr60 node_3 netRa60 -605178.5218201319
Lbr60 netRa60 netL60 9.265094484395861e-10
Rbbr60 netL60 0 2845420.5676623136
Cbr60 netL60 0 5.379670511670412e-22

* Branch 61
Rabr61 node_3 netRa61 2642109.450437911
Lbr61 netRa61 netL61 3.091439640407698e-09
Rbbr61 netL61 0 -4153493.415521572
Cbr61 netL61 0 2.8173776493542474e-22

* Branch 62
Rabr62 node_3 netRa62 1136602.596939116
Lbr62 netRa62 netL62 2.2639817171703633e-09
Rbbr62 netL62 0 -3127190.012282456
Cbr62 netL62 0 6.370723389464999e-22

* Branch 63
Rabr63 node_3 netRa63 -637224.6384791768
Lbr63 netRa63 netL63 1.158155060841128e-09
Rbbr63 netL63 0 3682572.7311121435
Cbr63 netL63 0 4.934647555229268e-22

* Branch 64
Rabr64 node_3 netRa64 -311088.8573712428
Lbr64 netRa64 netL64 1.1124888964708221e-09
Rbbr64 netL64 0 4774086.334706307
Cbr64 netL64 0 7.488500658579555e-22

* Branch 65
Rabr65 node_3 netRa65 -197999.35681966384
Lbr65 netRa65 netL65 1.0014879065768495e-09
Rbbr65 netL65 0 6472523.348002936
Cbr65 netL65 0 7.811527380487304e-22

* Branch 66
Rabr66 node_3 netRa66 -4909477.453370222
Lbr66 netRa66 netL66 1.4282513696816374e-09
Rbbr66 netL66 0 5900102.978005976
Cbr66 netL66 0 4.930602120818278e-23

* Branch 67
Rabr67 node_3 netRa67 -314539.6581751426
Lbr67 netRa67 netL67 1.358944161701918e-09
Rbbr67 netL67 0 6678687.4910151865
Cbr67 netL67 0 6.466823177442398e-22

* Branch 68
Rabr68 node_3 netRa68 4872054.323566128
Lbr68 netRa68 netL68 -1.9708454876688454e-09
Rbbr68 netL68 0 -6435389.804976946
Cbr68 netL68 0 -6.285701948415087e-23

* Branch 69
Rabr69 node_3 netRa69 -615585.3190767255
Lbr69 netRa69 netL69 1.438720276499478e-09
Rbbr69 netL69 0 6233007.69373386
Cbr69 netL69 0 3.749127435059239e-22

* Branch 70
Rabr70 node_3 netRa70 -5980202.060129148
Lbr70 netRa70 netL70 1.8275480083703454e-09
Rbbr70 netL70 0 7190702.198565121
Cbr70 netL70 0 4.2498577995626864e-23

* Branch 71
Rabr71 node_3 netRa71 -1690739.653546295
Lbr71 netRa71 netL71 -2.7699403976191384e-10
Rbbr71 netL71 0 1842482.1623564751
Cbr71 netL71 0 -8.891877866303592e-23

* Branch 72
Rabr72 node_3 netRa72 -451807.93869040336
Lbr72 netRa72 netL72 1.6323631855037374e-09
Rbbr72 netL72 0 10579643.68339402
Cbr72 netL72 0 3.414506890158613e-22

* Branch 73
Rabr73 node_3 netRa73 4678265853.061622
Lbr73 netRa73 netL73 -1.1290630887711176e-07
Rbbr73 netL73 0 -4679534176.272235
Cbr73 netL73 0 -5.157393784215e-27

* Branch 74
Rabr74 node_3 netRa74 526793.2192439277
Lbr74 netRa74 netL74 9.254973726536346e-10
Rbbr74 netL74 0 -2673958.2664064732
Cbr74 netL74 0 6.570647824306947e-22

* Branch 75
Rabr75 node_3 netRa75 -25465347.352018345
Lbr75 netRa75 netL75 4.4530230647357695e-09
Rbbr75 netL75 0 27112068.891013104
Cbr75 netL75 0 6.449706486029958e-24

* Branch 76
Rabr76 node_3 netRa76 92051.22809104683
Lbr76 netRa76 netL76 9.690088338876373e-10
Rbbr76 netL76 0 -10780124.174082952
Cbr76 netL76 0 9.768563398497405e-22

* Branch 77
Rabr77 node_3 netRa77 195101.17007428253
Lbr77 netRa77 netL77 1.1386780097701123e-09
Rbbr77 netL77 0 -8167175.333965012
Cbr77 netL77 0 7.146951415382158e-22

* Branch 78
Rabr78 node_3 netRa78 378297.59754482977
Lbr78 netRa78 netL78 8.985661701827393e-10
Rbbr78 netL78 0 -2855545.854718922
Cbr78 netL78 0 8.318489952757e-22

* Branch 79
Rabr79 node_3 netRa79 368208.25345628796
Lbr79 netRa79 netL79 2.214899390764458e-09
Rbbr79 netL79 0 -17411747.023611322
Cbr79 netL79 0 3.4548709751689787e-22

* Branch 80
Rabr80 node_3 netRa80 690097.5174015006
Lbr80 netRa80 netL80 9.226521646807452e-10
Rbbr80 netL80 0 -2370302.7624896783
Cbr80 netL80 0 5.640610903044929e-22

* Branch 81
Rabr81 node_3 netRa81 63319682.76458426
Lbr81 netRa81 netL81 5.449393617635319e-09
Rbbr81 netL81 0 -64361090.48902959
Cbr81 netL81 0 1.3371685056315156e-24

* Branch 82
Rabr82 node_3 netRa82 598571464.3740649
Lbr82 netRa82 netL82 -2.0059179393413626e-08
Rbbr82 netL82 0 -599958163.201586
Cbr82 netL82 0 -5.585681645574801e-26

* Branch 83
Rabr83 node_3 netRa83 -39957553.36924296
Lbr83 netRa83 netL83 2.281324964338328e-08
Rbbr83 netL83 0 45099927.3730204
Cbr83 netL83 0 1.2659370721443419e-23

* Branch 84
Rabr84 node_3 netRa84 614085734.0455116
Lbr84 netRa84 netL84 1.8036812701840953e-08
Rbbr84 netL84 0 -615290593.2308782
Cbr84 netL84 0 4.7736501017837485e-26

* Branch 85
Rabr85 node_3 netRa85 -44931422.22842339
Lbr85 netRa85 netL85 -8.68535843814187e-09
Rbbr85 netL85 0 48308544.413288176
Cbr85 netL85 0 -4.001423439492357e-24

* Branch 86
Rabr86 node_3 netRa86 324849.9203114443
Lbr86 netRa86 netL86 1.0221823714657186e-09
Rbbr86 netL86 0 -3576680.2214912027
Cbr86 netL86 0 8.797949400413963e-22

* Branch 87
Rabr87 node_3 netRa87 905771.592104359
Lbr87 netRa87 netL87 1.2678672930404432e-09
Rbbr87 netL87 0 -2636496.0304323626
Cbr87 netL87 0 5.30946834846941e-22

* Branch 88
Rabr88 node_3 netRa88 59033246.41745451
Lbr88 netRa88 netL88 2.854239426938138e-09
Rbbr88 netL88 0 -59469311.96850658
Cbr88 netL88 0 8.13021203972001e-25

* Branch 89
Rabr89 node_3 netRa89 718238.5104779394
Lbr89 netRa89 netL89 -1.1687780595561425e-09
Rbbr89 netL89 0 -4166016.6187889413
Cbr89 netL89 0 -3.9057266236420586e-22

* Branch 90
Rabr90 node_3 netRa90 13426921.542019265
Lbr90 netRa90 netL90 -3.4998128020128458e-09
Rbbr90 netL90 0 -14909164.273858426
Cbr90 netL90 0 -1.7482680816929884e-23

* Branch 91
Rabr91 node_3 netRa91 1775482.3149229793
Lbr91 netRa91 netL91 1.5449244756872393e-09
Rbbr91 netL91 0 -3039260.811859125
Cbr91 netL91 0 2.863169289630823e-22

* Branch 92
Rabr92 node_3 netRa92 469019.86683300586
Lbr92 netRa92 netL92 -1.3352836022729818e-09
Rbbr92 netL92 0 -7177153.048887971
Cbr92 netL92 0 -3.9659511068215245e-22

* Branch 93
Rabr93 node_3 netRa93 3545827.7538706725
Lbr93 netRa93 netL93 -2.0189039180044626e-09
Rbbr93 netL93 0 -5259083.344659603
Cbr93 netL93 0 -1.0826035853717505e-22

* Branch 94
Rabr94 node_3 netRa94 -10429561.345419643
Lbr94 netRa94 netL94 1.2626452405668481e-09
Rbbr94 netL94 0 10884130.52372111
Cbr94 netL94 0 1.1122783970435996e-23

* Branch 95
Rabr95 node_3 netRa95 299665.5220729795
Lbr95 netRa95 netL95 -3.0506464715236944e-10
Rbbr95 netL95 0 -1128428.8158563352
Cbr95 netL95 0 -9.018950315256381e-22

* Branch 96
Rabr96 node_3 netRa96 -20265467.526718497
Lbr96 netRa96 netL96 -1.0033644978881505e-09
Rbbr96 netL96 0 20387002.99635025
Cbr96 netL96 0 -2.4285963624193332e-24

* Branch 97
Rabr97 node_3 netRa97 -557913.0921068708
Lbr97 netRa97 netL97 -7.810460688714177e-10
Rbbr97 netL97 0 3350500.880251797
Cbr97 netL97 0 -4.1804825539775066e-22

* Branch 98
Rabr98 node_3 netRa98 124643.82440573045
Lbr98 netRa98 netL98 -2.698672933414127e-10
Rbbr98 netL98 0 -1717275.5927845899
Cbr98 netL98 0 -1.2594594134017133e-21

* Branch 99
Rabr99 node_3 netRa99 2262556.451342034
Lbr99 netRa99 netL99 1.700424121144635e-10
Rbbr99 netL99 0 -2307655.191046777
Cbr99 netL99 0 3.257718152839554e-23

.ends


* Y'34
.subckt yp34 node_3 node_4
* Branch 0
Rabr0 node_3 netRa0 -422.2397401554033
Lbr0 netRa0 netL0 2.0449866647844864e-13
Rbbr0 netL0 node_4 581.23871531924
Cbr0 netL0 node_4 7.767476697579449e-19

* Branch 1
Rabr1 node_3 netRa1 -1796.9804501316326
Lbr1 netRa1 netL1 3.6898914830691153e-13
Rbbr1 netL1 node_4 1924.764257518875
Cbr1 netL1 node_4 1.0381739811955911e-19

* Branch 2
Rabr2 node_3 netRa2 -374.04441088361597
Lbr2 netRa2 netL2 -2.613907947387005e-13
Rbbr2 netL2 node_4 732.9689471083525
Cbr2 netL2 node_4 -1.0398917788508737e-18

* Branch 3
Rabr3 node_3 netRa3 -19.45887224988599
Lbr3 netRa3 netL3 -2.1828865427068294e-13
Rbbr3 netL3 node_4 -28869.973853092346
Cbr3 netL3 node_4 -2.508574738346214e-18

* Branch 4
Rabr4 node_3 netRa4 -53.706618493769284
Lbr4 netRa4 netL4 -1.1096522523641395e-13
Rbbr4 netL4 node_4 564.0311832817906
Cbr4 netL4 node_4 -4.541919555594779e-18

* Branch 5
Rabr5 node_3 netRa5 -114.73418496010777
Lbr5 netRa5 netL5 -8.352253324756213e-14
Rbbr5 netL5 node_4 229.20970994775325
Cbr5 netL5 node_4 -3.3980553022043302e-18

* Branch 6
Rabr6 node_3 netRa6 65.821754941753
Lbr6 netRa6 netL6 -7.060595238247276e-14
Rbbr6 netL6 node_4 -194.69928801832236
Cbr6 netL6 node_4 -5.192034675866841e-18

* Branch 7
Rabr7 node_3 netRa7 99.48748804099162
Lbr7 netRa7 netL7 -6.405221866662686e-14
Rbbr7 netL7 node_4 -163.58361781923492
Cbr7 netL7 node_4 -3.826319667630178e-18

* Branch 8
Rabr8 node_3 netRa8 49.913655076632814
Lbr8 netRa8 netL8 6.21736685307915e-14
Rbbr8 netL8 node_4 -175.12044762530925
Cbr8 netL8 node_4 7.48288580850201e-18

* Branch 9
Rabr9 node_3 netRa9 71.62752830348103
Lbr9 netRa9 netL9 9.18388100642186e-14
Rbbr9 netL9 node_4 -266.9176581172282
Cbr9 netL9 node_4 5.0578722435161295e-18

* Branch 10
Rabr10 node_3 netRa10 -383.83289076326696
Lbr10 netRa10 netL10 1.164353270421218e-13
Rbbr10 netL10 node_4 439.4079685526779
Cbr10 netL10 node_4 6.834554840406329e-19

* Branch 11
Rabr11 node_3 netRa11 146.82894575491494
Lbr11 netRa11 netL11 1.5244518973179587e-13
Rbbr11 netL11 node_4 -429.5561278098801
Cbr11 netL11 node_4 2.5008867511434114e-18

* Branch 12
Rabr12 node_3 netRa12 9628.628553664024
Lbr12 netRa12 netL12 7.852220122555816e-13
Rbbr12 netL12 node_4 -9729.209316960338
Cbr12 netL12 node_4 8.401267613584405e-21

* Branch 13
Rabr13 node_3 netRa13 -33.46066525434657
Lbr13 netRa13 netL13 8.543079631639305e-14
Rbbr13 netL13 node_4 400.4718683708397
Cbr13 netL13 node_4 5.978266850428422e-18

* Branch 14
Rabr14 node_3 netRa14 -137.62718571869448
Lbr14 netRa14 netL14 -4.265013132726897e-13
Rbbr14 netL14 node_4 2181.485343803979
Cbr14 netL14 node_4 -1.542111005434939e-18

* Branch 15
Rabr15 node_3 netRa15 -14.091263835134933
Lbr15 netRa15 netL15 4.83521259388662e-14
Rbbr15 netL15 node_4 296.72164538744477
Cbr15 netL15 node_4 1.064156563299078e-17

* Branch 16
Rabr16 node_3 netRa16 -114.26004006946934
Lbr16 netRa16 netL16 -6.973323095521158e-14
Rbbr16 netL16 node_4 181.59006375082615
Cbr16 netL16 node_4 -3.407326357255027e-18

* Branch 17
Rabr17 node_3 netRa17 -2757.24530778853
Lbr17 netRa17 netL17 1.453107431396411e-12
Rbbr17 netL17 node_4 5067.414720361193
Cbr17 netL17 node_4 1.0283076206703223e-19

* Branch 18
Rabr18 node_3 netRa18 -105.11327545899616
Lbr18 netRa18 netL18 2.4593445914011397e-13
Rbbr18 netL18 node_4 1820.404208636927
Cbr18 netL18 node_4 1.2240590660075122e-18

* Branch 19
Rabr19 node_3 netRa19 -2224.9107211860987
Lbr19 netRa19 netL19 -1.2734939311445804e-12
Rbbr19 netL19 node_4 3226.4128794598555
Cbr19 netL19 node_4 -1.7959978035357357e-19

* Branch 20
Rabr20 node_3 netRa20 6112.543721678878
Lbr20 netRa20 netL20 -1.1736060332213782e-12
Rbbr20 netL20 node_4 -6862.075665506314
Cbr20 netL20 node_4 -2.7869939734712134e-20

* Branch 21
Rabr21 node_3 netRa21 -102.07851820179269
Lbr21 netRa21 netL21 -1.0498450579898972e-13
Rbbr21 netL21 node_4 269.4135277111618
Cbr21 netL21 node_4 -3.895638432504231e-18

* Branch 22
Rabr22 node_3 netRa22 -694.24007719261
Lbr22 netRa22 netL22 9.507359481166022e-13
Rbbr22 netL22 node_4 4769.7227870745555
Cbr22 netL22 node_4 2.7967550338422403e-19

* Branch 23
Rabr23 node_3 netRa23 -3105.838681006386
Lbr23 netRa23 netL23 -1.4906912874782056e-12
Rbbr23 netL23 node_4 5258.093128758982
Cbr23 netL23 node_4 -9.212828603731638e-20

* Branch 24
Rabr24 node_3 netRa24 -73.90167858875023
Lbr24 netRa24 netL24 -2.5177379412397153e-13
Rbbr24 netL24 node_4 1427.7229754287343
Cbr24 netL24 node_4 -2.5447395204428866e-18

* Branch 25
Rabr25 node_3 netRa25 -4958.635552694837
Lbr25 netRa25 netL25 -1.7307959766689243e-12
Rbbr25 netL25 node_4 6728.251414501502
Cbr25 netL25 node_4 -5.2192928053021163e-20

* Branch 26
Rabr26 node_3 netRa26 13030.575433402431
Lbr26 netRa26 netL26 1.7158728770713415e-12
Rbbr26 netL26 node_4 -13773.890817823862
Cbr26 netL26 node_4 9.581129807047798e-21

* Branch 27
Rabr27 node_3 netRa27 114.80067510503466
Lbr27 netRa27 netL27 6.600332014612686e-14
Rbbr27 netL27 node_4 -187.37460627944037
Cbr27 netL27 node_4 3.0969166216660495e-18

* Branch 28
Rabr28 node_3 netRa28 56608.16526959259
Lbr28 netRa28 netL28 -4.616565561605824e-12
Rbbr28 netL28 node_4 -57896.31742761302
Cbr28 netL28 node_4 -1.4068955854710042e-21

* Branch 29
Rabr29 node_3 netRa29 -494.9115341399517
Lbr29 netRa29 netL29 3.2803891251200145e-13
Rbbr29 netL29 node_4 987.566545406244
Cbr29 netL29 node_4 6.646105367201511e-19

* Branch 30
Rabr30 node_3 netRa30 -3232.030871517594
Lbr30 netRa30 netL30 -1.0436028098055292e-12
Rbbr30 netL30 node_4 3671.9458302492158
Cbr30 netL30 node_4 -8.835771724159452e-20

* Branch 31
Rabr31 node_3 netRa31 19609.873878583552
Lbr31 netRa31 netL31 -1.2923299982193058e-11
Rbbr31 netL31 node_4 -23521.42291934754
Cbr31 netL31 node_4 -2.777464487786636e-20

* Branch 32
Rabr32 node_3 netRa32 1425.6552734429188
Lbr32 netRa32 netL32 5.635057099365315e-13
Rbbr32 netL32 node_4 -1984.8978741230471
Cbr32 netL32 node_4 2.0014378026315723e-19

* Branch 33
Rabr33 node_3 netRa33 -1708.0946245620091
Lbr33 netRa33 netL33 7.813919457855307e-13
Rbbr33 netL33 node_4 2635.4516357120187
Cbr33 netL33 node_4 1.725836246175099e-19

* Branch 34
Rabr34 node_3 netRa34 -74.65923076495194
Lbr34 netRa34 netL34 -1.023918449797307e-12
Rbbr34 netL34 node_4 14357.857451391517
Cbr34 netL34 node_4 -1.1528753495689418e-18

* Branch 35
Rabr35 node_3 netRa35 -76.86844540626505
Lbr35 netRa35 netL35 1.2961568755026616e-13
Rbbr35 netL35 node_4 533.9618543102304
Cbr35 netL35 node_4 3.099208838667937e-18

* Branch 36
Rabr36 node_3 netRa36 2333.194608600065
Lbr36 netRa36 netL36 -8.833056605456715e-13
Rbbr36 netL36 node_4 -3313.3187304973994
Cbr36 netL36 node_4 -1.137863652318316e-19

* Branch 37
Rabr37 node_3 netRa37 101328.20248154666
Lbr37 netRa37 netL37 4.9946499036383235e-12
Rbbr37 netL37 node_4 -102106.34154455831
Cbr37 netL37 node_4 4.830065936712253e-22

* Branch 38
Rabr38 node_3 netRa38 10873.4778814897
Lbr38 netRa38 netL38 1.4106550500420133e-12
Rbbr38 netL38 node_4 -11318.865166518894
Cbr38 netL38 node_4 1.1476392668071898e-20

* Branch 39
Rabr39 node_3 netRa39 15658.665730713763
Lbr39 netRa39 netL39 -2.2310090659846975e-12
Rbbr39 netL39 node_4 -16680.126184228542
Cbr39 netL39 node_4 -8.529963222188997e-21

* Branch 40
Rabr40 node_3 netRa40 166.74349653332496
Lbr40 netRa40 netL40 -1.7303169628087047e-13
Rbbr40 netL40 node_4 -385.20442232954065
Cbr40 netL40 node_4 -2.6678421176348847e-18

* Branch 41
Rabr41 node_3 netRa41 -288.3603119769122
Lbr41 netRa41 netL41 1.622265623604592e-13
Rbbr41 netL41 node_4 476.7159955794392
Cbr41 netL41 node_4 1.1739228691991573e-18

* Branch 42
Rabr42 node_3 netRa42 24.408347205104118
Lbr42 netRa42 netL42 -4.3551177272324574e-13
Rbbr42 netL42 node_4 -6751.735919394525
Cbr42 netL42 node_4 -2.2644083957003034e-18

* Branch 43
Rabr43 node_3 netRa43 -7.184680880991926
Lbr43 netRa43 netL43 1.0388644192657405e-13
Rbbr43 netL43 node_4 2910.7208573304088
Cbr43 netL43 node_4 4.393112954089434e-18

* Branch 44
Rabr44 node_3 netRa44 1669.7198927497843
Lbr44 netRa44 netL44 8.170714148441208e-13
Rbbr44 netL44 node_4 -2739.1194222842637
Cbr44 netL44 node_4 1.794025413521666e-19

* Branch 45
Rabr45 node_3 netRa45 150.1941762933588
Lbr45 netRa45 netL45 -1.1063346719522629e-13
Rbbr45 netL45 node_4 -305.6877488266278
Cbr45 netL45 node_4 -2.3959116179748435e-18

* Branch 46
Rabr46 node_3 netRa46 110624889.39372595
Lbr46 netRa46 netL46 1.8018753988343084e-10
Rbbr46 netL46 node_4 -110625638.47608984
Cbr46 netL46 node_4 1.47238570471569e-26

* Branch 47
Rabr47 node_3 netRa47 -541.8246233083732
Lbr47 netRa47 netL47 3.102006849209523e-13
Rbbr47 netL47 node_4 955.0677915933219
Cbr47 netL47 node_4 5.971619649675417e-19

* Branch 48
Rabr48 node_3 netRa48 -24.001527671389397
Lbr48 netRa48 netL48 -1.5228501096668836e-12
Rbbr48 netL48 node_4 123242.510252488
Cbr48 netL48 node_4 -8.807477990912148e-19

* Branch 49
Rabr49 node_3 netRa49 -41.869130890951105
Lbr49 netRa49 netL49 -5.803591583416933e-13
Rbbr49 netL49 node_4 8087.934036853891
Cbr49 netL49 node_4 -1.8843924351378314e-18

* Branch 50
Rabr50 node_3 netRa50 43825.38464822381
Lbr50 netRa50 netL50 4.8926384837196234e-12
Rbbr50 netL50 node_4 -45735.37933423775
Cbr50 netL50 node_4 2.4427434565461822e-21

* Branch 51
Rabr51 node_3 netRa51 -107.04836087461914
Lbr51 netRa51 netL51 -2.4809874070466415e-13
Rbbr51 netL51 node_4 788.4536258371405
Cbr51 netL51 node_4 -2.983640839356214e-18

* Branch 52
Rabr52 node_3 netRa52 1281.8537244733975
Lbr52 netRa52 netL52 4.4767325985334866e-13
Rbbr52 netL52 node_4 -1630.1971119309965
Cbr52 netL52 node_4 2.1468404727768746e-19

* Branch 53
Rabr53 node_3 netRa53 43709.02618504695
Lbr53 netRa53 netL53 3.4178793382765105e-12
Rbbr53 netL53 node_4 -44018.85949981992
Cbr53 netL53 node_4 1.7771979979095272e-21

* Branch 54
Rabr54 node_3 netRa54 3346.6669949381367
Lbr54 netRa54 netL54 -1.0541393286589206e-12
Rbbr54 netL54 node_4 -4266.573915859343
Cbr54 netL54 node_4 -7.369947505576759e-20

* Branch 55
Rabr55 node_3 netRa55 2375.455170067534
Lbr55 netRa55 netL55 -9.97514844440708e-13
Rbbr55 netL55 node_4 -3560.6468917789475
Cbr55 netL55 node_4 -1.1766909347141142e-19

* Branch 56
Rabr56 node_3 netRa56 194.80278528668634
Lbr56 netRa56 netL56 -2.6940356736462325e-12
Rbbr56 netL56 node_4 -23796.587466191606
Cbr56 netL56 node_4 -5.423822182824463e-19

* Branch 57
Rabr57 node_3 netRa57 3919.06275670235
Lbr57 netRa57 netL57 -6.4089003684465135e-12
Rbbr57 netL57 node_4 -9657.136073569774
Cbr57 netL57 node_4 -1.680650722502695e-19

* Branch 58
Rabr58 node_3 netRa58 143.63115188055926
Lbr58 netRa58 netL58 -4.788610644922012e-13
Rbbr58 netL58 node_4 -4317.623035758778
Cbr58 netL58 node_4 -7.606191944677395e-19

* Branch 59
Rabr59 node_3 netRa59 1011987.6888480824
Lbr59 netRa59 netL59 -1.3260347025445744e-11
Rbbr59 netL59 node_4 -1012400.368696657
Cbr59 netL59 node_4 -1.294206739826632e-23

* Branch 60
Rabr60 node_3 netRa60 -12482.105960483954
Lbr60 netRa60 netL60 -2.464772689459708e-12
Rbbr60 netL60 node_4 13085.779875279584
Cbr60 netL60 node_4 -1.510097492366345e-20

* Branch 61
Rabr61 node_3 netRa61 10353.074409690042
Lbr61 netRa61 netL61 -3.832492967658702e-12
Rbbr61 netL61 node_4 -11938.993012014394
Cbr61 netL61 node_4 -3.097033687130011e-20

* Branch 62
Rabr62 node_3 netRa62 2028.2319559019586
Lbr62 netRa62 netL62 -9.769090604430102e-13
Rbbr62 netL62 node_4 -3305.9133738967453
Cbr62 netL62 node_4 -1.4548304433031923e-19

* Branch 63
Rabr63 node_3 netRa63 5179.437641089011
Lbr63 netRa63 netL63 2.174557125061494e-12
Rbbr63 netL63 node_4 -8433.983582655044
Cbr63 netL63 node_4 4.982754317291329e-20

* Branch 64
Rabr64 node_3 netRa64 2280.766535155978
Lbr64 netRa64 netL64 -1.1720637003804593e-12
Rbbr64 netL64 node_4 -3849.2442257357375
Cbr64 netL64 node_4 -1.3335016794179544e-19

* Branch 65
Rabr65 node_3 netRa65 1259.9598143569647
Lbr65 netRa65 netL65 -8.04864863884757e-13
Rbbr65 netL65 node_4 -2747.6635281080908
Cbr65 netL65 node_4 -2.322032437362376e-19

* Branch 66
Rabr66 node_3 netRa66 78837.57482635565
Lbr66 netRa66 netL66 2.397432542308969e-11
Rbbr66 netL66 node_4 -84486.03197205036
Cbr66 netL66 node_4 3.6014217631237265e-21

* Branch 67
Rabr67 node_3 netRa67 33.3965387788549
Lbr67 netRa67 netL67 -3.3008528433328126e-13
Rbbr67 netL67 node_4 -7485.54103726571
Cbr67 netL67 node_4 -1.2993536187104683e-18

* Branch 68
Rabr68 node_3 netRa68 137.33986620996285
Lbr68 netRa68 netL68 -4.413154054003245e-13
Rbbr68 netL68 node_4 -3339.155615457713
Cbr68 netL68 node_4 -9.576454987929987e-19

* Branch 69
Rabr69 node_3 netRa69 -1881.0570418428492
Lbr69 netRa69 netL69 -6.697052923513147e-13
Rbbr69 netL69 node_4 2347.4973408285655
Cbr69 netL69 node_4 -1.517378527515492e-19

* Branch 70
Rabr70 node_3 netRa70 13741.501543406572
Lbr70 netRa70 netL70 9.3929141658972e-12
Rbbr70 netL70 node_4 -18925.246633961626
Cbr70 netL70 node_4 3.61520465497652e-20

* Branch 71
Rabr71 node_3 netRa71 5102.402193594594
Lbr71 netRa71 netL71 9.167072376355607e-12
Rbbr71 netL71 node_4 -20635.381574082232
Cbr71 netL71 node_4 8.72623541230099e-20

* Branch 72
Rabr72 node_3 netRa72 1166.2380125099628
Lbr72 netRa72 netL72 -4.8824808818985014e-12
Rbbr72 netL72 node_4 -13244.69003189174
Cbr72 netL72 node_4 -3.1445912618097867e-19

* Branch 73
Rabr73 node_3 netRa73 2980.6789668708934
Lbr73 netRa73 netL73 3.645531611638602e-12
Rbbr73 netL73 node_4 -7492.080848966159
Cbr73 netL73 node_4 1.6348971187083667e-19

* Branch 74
Rabr74 node_3 netRa74 9452.881946328598
Lbr74 netRa74 netL74 1.0495395905920499e-11
Rbbr74 netL74 node_4 -21679.55390032165
Cbr74 netL74 node_4 5.1280118360496183e-20

* Branch 75
Rabr75 node_3 netRa75 983274.3505261623
Lbr75 netRa75 netL75 -7.893543325060125e-11
Rbbr75 netL75 node_4 -990142.0169826641
Cbr75 netL75 node_4 -8.1070311331095e-23

* Branch 76
Rabr76 node_3 netRa76 10897.583180961443
Lbr76 netRa76 netL76 -1.0817043343738298e-11
Rbbr76 netL76 node_4 -17585.824550440204
Cbr76 netL76 node_4 -5.6386591446959e-20

* Branch 77
Rabr77 node_3 netRa77 27921.24799559781
Lbr77 netRa77 netL77 -1.1968615237605378e-11
Rbbr77 netL77 node_4 -32216.637318098827
Cbr77 netL77 node_4 -1.3299624954213235e-20

* Branch 78
Rabr78 node_3 netRa78 1568.9554774647397
Lbr78 netRa78 netL78 5.4100226717794134e-12
Rbbr78 netL78 node_4 -24024.68811193928
Cbr78 netL78 node_4 1.4399723785425358e-19

* Branch 79
Rabr79 node_3 netRa79 5869.303267888444
Lbr79 netRa79 netL79 7.248688000925397e-12
Rbbr79 netL79 node_4 -14614.427545350778
Cbr79 netL79 node_4 8.460558472633138e-20

* Branch 80
Rabr80 node_3 netRa80 1672.955880027881
Lbr80 netRa80 netL80 -5.1320977861615425e-12
Rbbr80 netL80 node_4 -10997.581178124952
Cbr80 netL80 node_4 -2.786005506792822e-19

* Branch 81
Rabr81 node_3 netRa81 17409.639537515854
Lbr81 netRa81 netL81 -1.6521458012568567e-11
Rbbr81 netL81 node_4 -31062.202683095024
Cbr81 netL81 node_4 -3.0540256979652213e-20

* Branch 82
Rabr82 node_3 netRa82 5930.655715124641
Lbr82 netRa82 netL82 -5.685701826294731e-12
Rbbr82 netL82 node_4 -10860.222722963592
Cbr82 netL82 node_4 -8.826033269585625e-20

* Branch 83
Rabr83 node_3 netRa83 2072.4887331761533
Lbr83 netRa83 netL83 -7.782293246667272e-12
Rbbr83 netL83 node_4 -22844.793594156676
Cbr83 netL83 node_4 -1.6427331118252946e-19

* Branch 84
Rabr84 node_3 netRa84 2050.768393831999
Lbr84 netRa84 netL84 -9.5155420902444e-12
Rbbr84 netL84 node_4 -30824.086974714915
Cbr84 netL84 node_4 -1.5043734606987538e-19

* Branch 85
Rabr85 node_3 netRa85 3235.650049090496
Lbr85 netRa85 netL85 -1.8829006390308092e-11
Rbbr85 netL85 node_4 -59677.116418688965
Cbr85 netL85 node_4 -9.747152432553939e-20

* Branch 86
Rabr86 node_3 netRa86 376.4408985360869
Lbr86 netRa86 netL86 -6.953791130911291e-12
Rbbr86 netL86 node_4 -53915.60012118112
Cbr86 netL86 node_4 -3.4241592627224454e-19

* Branch 87
Rabr87 node_3 netRa87 431.37948885828297
Lbr87 netRa87 netL87 -5.724181017957198e-12
Rbbr87 netL87 node_4 -37585.824937147714
Cbr87 netL87 node_4 -3.5289560831295163e-19

* Branch 88
Rabr88 node_3 netRa88 499.14500448663347
Lbr88 netRa88 netL88 -6.045934148172802e-12
Rbbr88 netL88 node_4 -32753.848051000914
Cbr88 netL88 node_4 -3.6974068381026173e-19

* Branch 89
Rabr89 node_3 netRa89 3843.79102627604
Lbr89 netRa89 netL89 -1.5609779840264548e-11
Rbbr89 netL89 node_4 -38159.48948209941
Cbr89 netL89 node_4 -1.0640333584812542e-19

* Branch 90
Rabr90 node_3 netRa90 2857.109250873134
Lbr90 netRa90 netL90 -6.237743761684562e-12
Rbbr90 netL90 node_4 -12125.700591428473
Cbr90 netL90 node_4 -1.8002356749548784e-19

* Branch 91
Rabr91 node_3 netRa91 478.5339310368719
Lbr91 netRa91 netL91 -3.5358368618231976e-12
Rbbr91 netL91 node_4 -12598.191136362504
Cbr91 netL91 node_4 -5.858098030212548e-19

* Branch 92
Rabr92 node_3 netRa92 1493.392896879871
Lbr92 netRa92 netL92 -2.8464576255488168e-12
Rbbr92 netL92 node_4 -5511.182019166581
Cbr92 netL92 node_4 -3.457407880289717e-19

* Branch 93
Rabr93 node_3 netRa93 2441.4548292378463
Lbr93 netRa93 netL93 -7.092440901996743e-12
Rbbr93 netL93 node_4 -14132.419245815383
Cbr93 netL93 node_4 -2.0545098738860999e-19

* Branch 94
Rabr94 node_3 netRa94 793.4872233075292
Lbr94 netRa94 netL94 2.7986303711808433e-12
Rbbr94 netL94 node_4 -4697.766571188798
Cbr94 netL94 node_4 7.52314219872499e-19

* Branch 95
Rabr95 node_3 netRa95 6662459.306447585
Lbr95 netRa95 netL95 -1.6457521499158134e-10
Rbbr95 netL95 node_4 -6667656.844981346
Cbr95 netL95 node_4 -3.7046755263074455e-24

* Branch 96
Rabr96 node_3 netRa96 -1372.4081037363258
Lbr96 netRa96 netL96 -6.192385270668888e-13
Rbbr96 netL96 node_4 1933.3301662540841
Cbr96 netL96 node_4 -2.3352535651013767e-19

* Branch 97
Rabr97 node_3 netRa97 -3365.5511545259783
Lbr97 netRa97 netL97 -4.535432343783569e-13
Rbbr97 netL97 node_4 3490.316997653781
Cbr97 netL97 node_4 -3.8616973342451486e-20

* Branch 98
Rabr98 node_3 netRa98 77.21950117202087
Lbr98 netRa98 netL98 7.504453780788112e-14
Rbbr98 netL98 node_4 -197.96332913508957
Cbr98 netL98 node_4 5.2142634326264925e-18

* Branch 99
Rabr99 node_3 netRa99 -1068.764890008296
Lbr99 netRa99 netL99 -2.5590609826171966e-13
Rbbr99 netL99 node_4 1178.9788929525114
Cbr99 netL99 node_4 -2.0859472793152073e-19

.ends


* Y'44
.subckt yp44 node_4 0
* Branch 0
Rabr0 node_4 netRa0 71963.36659575586
Lbr0 netRa0 netL0 -5.532867435088293e-11
Rbbr0 netL0 0 -203831.96656265337
Cbr0 netL0 0 -3.7044636681814384e-21

* Branch 1
Rabr1 node_4 netRa1 2111724.033559289
Lbr1 netRa1 netL1 -2.4021384920701294e-10
Rbbr1 netL1 0 -2179196.263369425
Cbr1 netL1 0 -5.2064845958500397e-23

* Branch 2
Rabr2 node_4 netRa2 53062.54709095622
Lbr2 netRa2 netL2 -5.3332310627255964e-11
Rbbr2 netL2 0 -171916.43760380472
Cbr2 netL2 0 -5.718313155890976e-21

* Branch 3
Rabr3 node_4 netRa3 25204.070772969913
Lbr3 netRa3 netL3 -3.4126214111322543e-11
Rbbr3 netL3 0 -140241.34825468462
Cbr3 netL3 0 -9.380310091691016e-21

* Branch 4
Rabr4 node_4 netRa4 69377.06354011122
Lbr4 netRa4 netL4 -5.214142026594747e-11
Rbbr4 netL4 0 -161635.1259680978
Cbr4 netL4 0 -4.577281661709766e-21

* Branch 5
Rabr5 node_4 netRa5 14208.37423875494
Lbr5 netRa5 netL5 -1.8245850282920563e-11
Rbbr5 netL5 0 -91593.6314673795
Cbr5 netL5 0 -1.3660684632294032e-20

* Branch 6
Rabr6 node_4 netRa6 16736398.599288713
Lbr6 netRa6 netL6 4.807967175477293e-10
Rbbr6 netL6 0 -16778360.81744376
Cbr6 netL6 0 1.7130468622717692e-24

* Branch 7
Rabr7 node_4 netRa7 22187.82843662754
Lbr7 netRa7 netL7 -6.377990450933926e-11
Rbbr7 netL7 0 -496139.5057397884
Cbr7 netL7 0 -5.534492004212897e-21

* Branch 8
Rabr8 node_4 netRa8 -31880.94289538875
Lbr8 netRa8 netL8 -1.1417263457683713e-10
Rbbr8 netL8 0 465779.88219655183
Cbr8 netL8 0 -8.16433085090411e-21

* Branch 9
Rabr9 node_4 netRa9 32224.43962923799
Lbr9 netRa9 netL9 -6.84880853436672e-11
Rbbr9 netL9 0 -306955.48707482603
Cbr9 netL9 0 -6.693397856216062e-21

* Branch 10
Rabr10 node_4 netRa10 30280.879272972074
Lbr10 netRa10 netL10 -2.7792730217225346e-11
Rbbr10 netL10 0 -104462.73777188582
Cbr10 netL10 0 -8.665919721662283e-21

* Branch 11
Rabr11 node_4 netRa11 -13069.62596551647
Lbr11 netRa11 netL11 -1.0019197873213806e-10
Rbbr11 netL11 0 1001331.0738017028
Cbr11 netL11 0 -8.657482095254183e-21

* Branch 12
Rabr12 node_4 netRa12 69286.56887276501
Lbr12 netRa12 netL12 -1.3666680568049695e-10
Rbbr12 netL12 0 -411463.44593906775
Cbr12 netL12 0 -4.660393558303535e-21

* Branch 13
Rabr13 node_4 netRa13 16062.43937126366
Lbr13 netRa13 netL13 -6.94218098490199e-11
Rbbr13 netL13 0 -347575.5654997362
Cbr13 netL13 0 -1.1704619817283746e-20

* Branch 14
Rabr14 node_4 netRa14 345423.2640074854
Lbr14 netRa14 netL14 2.4837278865559634e-10
Rbbr14 netL14 0 -514781.26408189186
Cbr14 netL14 0 1.4109011821051706e-21

* Branch 15
Rabr15 node_4 netRa15 56888.19975729465
Lbr15 netRa15 netL15 4.1512907286122315e-11
Rbbr15 netL15 0 -137271.1111232673
Cbr15 netL15 0 5.368912179079882e-21

* Branch 16
Rabr16 node_4 netRa16 29793.884807961174
Lbr16 netRa16 netL16 -1.1026090135594728e-10
Rbbr16 netL16 0 -352102.10604343255
Cbr16 netL16 0 -1.0026616356543828e-20

* Branch 17
Rabr17 node_4 netRa17 13144.035107226604
Lbr17 netRa17 netL17 -1.0425772397268142e-10
Rbbr17 netL17 0 -816817.6045853934
Cbr17 netL17 0 -8.808215822475084e-21

* Branch 18
Rabr18 node_4 netRa18 -371139.35057282884
Lbr18 netRa18 netL18 -2.3032626050155079e-10
Rbbr18 netL18 0 510430.2468579629
Cbr18 netL18 0 -1.2256433352651938e-21

* Branch 19
Rabr19 node_4 netRa19 52670.95162109804
Lbr19 netRa19 netL19 -1.1132406167174898e-10
Rbbr19 netL19 0 -256321.51341823835
Cbr19 netL19 0 -8.028825915694953e-21

* Branch 20
Rabr20 node_4 netRa20 31658.854181627354
Lbr20 netRa20 netL20 -6.81179927620284e-11
Rbbr20 netL20 0 -291688.0525961622
Cbr20 netL20 0 -7.180435966766195e-21

* Branch 21
Rabr21 node_4 netRa21 19369.554294343667
Lbr21 netRa21 netL21 -2.4904618737112398e-11
Rbbr21 netL21 0 -115917.84836091347
Cbr21 netL21 0 -1.0917369141891508e-20

* Branch 22
Rabr22 node_4 netRa22 32288.678974286886
Lbr22 netRa22 netL22 -1.3123031125394194e-10
Rbbr22 netL22 0 -374024.8367979158
Cbr22 netL22 0 -1.0352262135242441e-20

* Branch 23
Rabr23 node_4 netRa23 21885.82007668188
Lbr23 netRa23 netL23 -7.874870232218407e-11
Rbbr23 netL23 0 -463817.24248506094
Cbr23 netL23 0 -7.431301857439546e-21

* Branch 24
Rabr24 node_4 netRa24 -143852.40816314926
Lbr24 netRa24 netL24 -1.6718407954747972e-10
Rbbr24 netL24 0 289295.7850286108
Cbr24 netL24 0 -4.073716801682964e-21

* Branch 25
Rabr25 node_4 netRa25 23965.49854134454
Lbr25 netRa25 netL25 -7.877393336111419e-11
Rbbr25 netL25 0 -404599.7763744217
Cbr25 netL25 0 -7.825941303750265e-21

* Branch 26
Rabr26 node_4 netRa26 -102335.92485919096
Lbr26 netRa26 netL26 -6.074748274872574e-11
Rbbr26 netL26 0 230098.306022793
Cbr26 netL26 0 -2.597581738087799e-21

* Branch 27
Rabr27 node_4 netRa27 -161257.44178786618
Lbr27 netRa27 netL27 -2.520854118615826e-10
Rbbr27 netL27 0 447506.871498677
Cbr27 netL27 0 -3.556873807092628e-21

* Branch 28
Rabr28 node_4 netRa28 11345.753668027142
Lbr28 netRa28 netL28 -1.5140506223334298e-10
Rbbr28 netL28 0 -982258.7237932401
Cbr28 netL28 0 -1.1850015383663856e-20

* Branch 29
Rabr29 node_4 netRa29 12698.588097170008
Lbr29 netRa29 netL29 -8.346394840318002e-11
Rbbr29 netL29 0 -747970.8697747713
Cbr29 netL29 0 -8.198567330106124e-21

* Branch 30
Rabr30 node_4 netRa30 61443.95255871822
Lbr30 netRa30 netL30 -8.11306167517812e-11
Rbbr30 netL30 0 -106052.26177408473
Cbr30 netL30 0 -1.228050648386086e-20

* Branch 31
Rabr31 node_4 netRa31 18034.262062934562
Lbr31 netRa31 netL31 -1.4804299384565613e-10
Rbbr31 netL31 0 -698461.832968582
Cbr31 netL31 0 -1.0826155247230261e-20

* Branch 32
Rabr32 node_4 netRa32 -826239.8894373976
Lbr32 netRa32 netL32 -8.313681121351438e-10
Rbbr32 netL32 0 1981182.2112138593
Cbr32 netL32 0 -5.127821894675539e-22

* Branch 33
Rabr33 node_4 netRa33 22788.03735785714
Lbr33 netRa33 netL33 -9.055190939639633e-11
Rbbr33 netL33 0 -291803.1711106348
Cbr33 netL33 0 -1.3153222055800121e-20

* Branch 34
Rabr34 node_4 netRa34 29612.431182733522
Lbr34 netRa34 netL34 -7.369973758082302e-11
Rbbr34 netL34 0 -339245.0532831207
Cbr34 netL34 0 -7.187533157220503e-21

* Branch 35
Rabr35 node_4 netRa35 34582.85818180287
Lbr35 netRa35 netL35 -5.903021349556485e-11
Rbbr35 netL35 0 -237825.66071321504
Cbr35 netL35 0 -7.084051360878792e-21

* Branch 36
Rabr36 node_4 netRa36 -16235.473350950986
Lbr36 netRa36 netL36 -7.502687618760943e-11
Rbbr36 netL36 0 380971.0446998983
Cbr36 netL36 0 -1.2548430962683347e-20

* Branch 37
Rabr37 node_4 netRa37 13854.00675171508
Lbr37 netRa37 netL37 -4.770259654529278e-11
Rbbr37 netL37 0 -457347.33154242206
Cbr37 netL37 0 -7.358655885623247e-21

* Branch 38
Rabr38 node_4 netRa38 29283.08441849873
Lbr38 netRa38 netL38 -8.063303574642834e-11
Rbbr38 netL38 0 -299796.59983324294
Cbr38 netL38 0 -9.027905538649127e-21

* Branch 39
Rabr39 node_4 netRa39 162824.1163356818
Lbr39 netRa39 netL39 -1.5741918376163442e-10
Rbbr39 netL39 0 -235232.49203588054
Cbr39 netL39 0 -4.085529951502078e-21

* Branch 40
Rabr40 node_4 netRa40 5755.804631887174
Lbr40 netRa40 netL40 -6.791722098710198e-11
Rbbr40 netL40 0 -575423.9899967099
Cbr40 netL40 0 -1.9175698214079385e-20

* Branch 41
Rabr41 node_4 netRa41 40223.81171157759
Lbr41 netRa41 netL41 -5.373706499837286e-11
Rbbr41 netL41 0 -196789.68344439403
Cbr41 netL41 0 -6.744641958373974e-21

* Branch 42
Rabr42 node_4 netRa42 9094.62521255127
Lbr42 netRa42 netL42 -1.18794911090893e-11
Rbbr42 netL42 0 -59329.0117813321
Cbr42 netL42 0 -2.1877857161061444e-20

* Branch 43
Rabr43 node_4 netRa43 22007.302300165124
Lbr43 netRa43 netL43 -2.0367600714624483e-11
Rbbr43 netL43 0 -83920.5484911531
Cbr43 netL43 0 -1.0984199657837842e-20

* Branch 44
Rabr44 node_4 netRa44 86048.82018574173
Lbr44 netRa44 netL44 -1.468492292525394e-10
Rbbr44 netL44 0 -286508.080210695
Cbr44 netL44 0 -5.9129481152301725e-21

* Branch 45
Rabr45 node_4 netRa45 241993.59552825996
Lbr45 netRa45 netL45 -1.9202890179377731e-10
Rbbr45 netL45 0 -345977.0089844576
Cbr45 netL45 0 -2.2858130902000642e-21

* Branch 46
Rabr46 node_4 netRa46 -5183.96789230015
Lbr46 netRa46 netL46 -1.2481930159346918e-10
Rbbr46 netL46 0 2176008.5718258508
Cbr46 netL46 0 -1.2281865763903893e-20

* Branch 47
Rabr47 node_4 netRa47 613501.9926156068
Lbr47 netRa47 netL47 -1.7629504250893763e-10
Rbbr47 netL47 0 -710092.9394505272
Cbr47 netL47 0 -4.042220827943098e-22

* Branch 48
Rabr48 node_4 netRa48 56549.23936340275
Lbr48 netRa48 netL48 -6.574453597897818e-11
Rbbr48 netL48 0 -158951.73571304444
Cbr48 netL48 0 -7.282631492952478e-21

* Branch 49
Rabr49 node_4 netRa49 -229407.178867061
Lbr49 netRa49 netL49 -1.6198492732583815e-10
Rbbr49 netL49 0 569414.1095937615
Cbr49 netL49 0 -1.2429387783083574e-21

* Branch 50
Rabr50 node_4 netRa50 27476.916527636837
Lbr50 netRa50 netL50 -1.1056684155828922e-10
Rbbr50 netL50 0 -222408.46742322657
Cbr50 netL50 0 -1.7856939775435272e-20

* Branch 51
Rabr51 node_4 netRa51 91940.37236448335
Lbr51 netRa51 netL51 9.415709006202496e-11
Rbbr51 netL51 0 -317293.5722879709
Cbr51 netL51 0 3.238236616989171e-21

* Branch 52
Rabr52 node_4 netRa52 47596.392011230295
Lbr52 netRa52 netL52 -4.20465829962359e-11
Rbbr52 netL52 0 -176830.57349623894
Cbr52 netL52 0 -4.981923613600557e-21

* Branch 53
Rabr53 node_4 netRa53 243631.78639503603
Lbr53 netRa53 netL53 -1.9258683774409165e-10
Rbbr53 netL53 0 -381385.21842528606
Cbr53 netL53 0 -2.0679943973498597e-21

* Branch 54
Rabr54 node_4 netRa54 161119.19025047673
Lbr54 netRa54 netL54 -1.1857971838603237e-10
Rbbr54 netL54 0 -373742.1186404921
Cbr54 netL54 0 -1.9655267295106427e-21

* Branch 55
Rabr55 node_4 netRa55 -105702.36572429925
Lbr55 netRa55 netL55 2.9109648147239545e-11
Rbbr55 netL55 0 133849.10436622016
Cbr55 netL55 0 2.0560721515842437e-21

* Branch 56
Rabr56 node_4 netRa56 2197767.6391141308
Lbr56 netRa56 netL56 3.827675102723776e-10
Rbbr56 netL56 0 -2387772.7547273487
Cbr56 netL56 0 7.296481790481566e-23

* Branch 57
Rabr57 node_4 netRa57 -257577.5423517053
Lbr57 netRa57 netL57 -2.960830028383796e-10
Rbbr57 netL57 0 428630.8791719713
Cbr57 netL57 0 -2.6870899022554663e-21

* Branch 58
Rabr58 node_4 netRa58 171856.76808795726
Lbr58 netRa58 netL58 -1.3858914213276672e-10
Rbbr58 netL58 0 -413851.08490109094
Cbr58 netL58 0 -1.9459050354125413e-21

* Branch 59
Rabr59 node_4 netRa59 -545913.2058130659
Lbr59 netRa59 netL59 -4.839550547765884e-10
Rbbr59 netL59 0 766774.6167870347
Cbr59 netL59 0 -1.1578895112846131e-21

* Branch 60
Rabr60 node_4 netRa60 67438.45129639923
Lbr60 netRa60 netL60 -1.2696656377594286e-10
Rbbr60 netL60 0 -635668.85521248
Cbr60 netL60 0 -2.9526803202464468e-21

* Branch 61
Rabr61 node_4 netRa61 -3918.550928562012
Lbr61 netRa61 netL61 -1.3766172455348793e-10
Rbbr61 netL61 0 14291089.369092472
Cbr61 netL61 0 -2.606834222332044e-21

* Branch 62
Rabr62 node_4 netRa62 152750.93801215437
Lbr62 netRa62 netL62 -1.8952944490640436e-10
Rbbr62 netL62 0 -513238.82008743647
Cbr62 netL62 0 -2.4134677536027308e-21

* Branch 63
Rabr63 node_4 netRa63 82152.44105439923
Lbr63 netRa63 netL63 -1.0255852708285505e-10
Rbbr63 netL63 0 -284487.1546160997
Cbr63 netL63 0 -4.380832760956068e-21

* Branch 64
Rabr64 node_4 netRa64 92251.6790801255
Lbr64 netRa64 netL64 -1.789883999479473e-10
Rbbr64 netL64 0 -578660.2067463106
Cbr64 netL64 0 -3.345598188566592e-21

* Branch 65
Rabr65 node_4 netRa65 61648.063871686536
Lbr65 netRa65 netL65 -1.2874801328425708e-10
Rbbr65 netL65 0 -343280.1339342991
Cbr65 netL65 0 -6.0697522029507746e-21

* Branch 66
Rabr66 node_4 netRa66 149341.24931576214
Lbr66 netRa66 netL66 -1.8433583556596965e-10
Rbbr66 netL66 0 -478305.1549817623
Cbr66 netL66 0 -2.5772814266115802e-21

* Branch 67
Rabr67 node_4 netRa67 62282.332039774374
Lbr67 netRa67 netL67 -2.43943914725763e-10
Rbbr67 netL67 0 -891887.887618032
Cbr67 netL67 0 -4.374570376148473e-21

* Branch 68
Rabr68 node_4 netRa68 180029.28893798558
Lbr68 netRa68 netL68 -1.667637898979032e-10
Rbbr68 netL68 0 -506467.3663527787
Cbr68 netL68 0 -1.827298851460318e-21

* Branch 69
Rabr69 node_4 netRa69 143684.71576081956
Lbr69 netRa69 netL69 -2.727282755739355e-10
Rbbr69 netL69 0 -577335.2182628851
Cbr69 netL69 0 -3.282992427000253e-21

* Branch 70
Rabr70 node_4 netRa70 109012.65651467013
Lbr70 netRa70 netL70 -1.453751589031897e-10
Rbbr70 netL70 0 -469587.7348229957
Cbr70 netL70 0 -2.8372631640014745e-21

* Branch 71
Rabr71 node_4 netRa71 -665307.8873800411
Lbr71 netRa71 netL71 -7.792977033934587e-10
Rbbr71 netL71 0 1159883.9187432108
Cbr71 netL71 0 -1.010536752264327e-21

* Branch 72
Rabr72 node_4 netRa72 197958.16885598731
Lbr72 netRa72 netL72 -2.1366691536356057e-10
Rbbr72 netL72 0 -661562.9101125814
Cbr72 netL72 0 -1.630546317870648e-21

* Branch 73
Rabr73 node_4 netRa73 131135.5223886483
Lbr73 netRa73 netL73 -1.7802370963629978e-10
Rbbr73 netL73 0 -534750.2188650002
Cbr73 netL73 0 -2.5368687789634132e-21

* Branch 74
Rabr74 node_4 netRa74 -147434.53837792855
Lbr74 netRa74 netL74 -4.715247913702724e-10
Rbbr74 netL74 0 1841791.1076975192
Cbr74 netL74 0 -1.7392322567458346e-21

* Branch 75
Rabr75 node_4 netRa75 -61293.658983545225
Lbr75 netRa75 netL75 -3.9300416863608914e-10
Rbbr75 netL75 0 1498088.0502246125
Cbr75 netL75 0 -4.292881335642334e-21

* Branch 76
Rabr76 node_4 netRa76 151025.66426742062
Lbr76 netRa76 netL76 -3.119301659728009e-10
Rbbr76 netL76 0 -849209.280821751
Cbr76 netL76 0 -2.4301951351142358e-21

* Branch 77
Rabr77 node_4 netRa77 -2750277.2026663767
Lbr77 netRa77 netL77 3.5893706662800023e-10
Rbbr77 netL77 0 2898441.3926099017
Cbr77 netL77 0 4.5025285749576663e-23

* Branch 78
Rabr78 node_4 netRa78 103684.0440635286
Lbr78 netRa78 netL78 -1.8506483108253438e-10
Rbbr78 netL78 0 -670703.3360440627
Cbr78 netL78 0 -2.6595235703755842e-21

* Branch 79
Rabr79 node_4 netRa79 -172858.27995475844
Lbr79 netRa79 netL79 -4.953601948647142e-10
Rbbr79 netL79 0 1019313.9774081169
Cbr79 netL79 0 -2.8142426185637064e-21

* Branch 80
Rabr80 node_4 netRa80 -271856.5981338499
Lbr80 netRa80 netL80 1.659963495038956e-10
Rbbr80 netL80 0 542478.43521282
Cbr80 netL80 0 1.1253403846224174e-21

* Branch 81
Rabr81 node_4 netRa81 -152515.51781950388
Lbr81 netRa81 netL81 -5.234346640309903e-10
Rbbr81 netL81 0 1273212.406691543
Cbr81 netL81 0 -2.697156774292704e-21

* Branch 82
Rabr82 node_4 netRa82 465198.9488173001
Lbr82 netRa82 netL82 -3.74012917077662e-10
Rbbr82 netL82 0 -849838.5694577477
Cbr82 netL82 0 -9.459964104763573e-22

* Branch 83
Rabr83 node_4 netRa83 62622.78169324881
Lbr83 netRa83 netL83 -8.644974377900451e-11
Rbbr83 netL83 0 -211055.4345167217
Cbr83 netL83 0 -6.540757267547185e-21

* Branch 84
Rabr84 node_4 netRa84 42397.51684447915
Lbr84 netRa84 netL84 -9.08146721823401e-11
Rbbr84 netL84 0 -276571.6983405735
Cbr84 netL84 0 -7.744258612392185e-21

* Branch 85
Rabr85 node_4 netRa85 53431.546217828356
Lbr85 netRa85 netL85 -1.3322536380372338e-10
Rbbr85 netL85 0 -184548.5094774517
Cbr85 netL85 0 -1.3508658598916173e-20

* Branch 86
Rabr86 node_4 netRa86 627901.6380936092
Lbr86 netRa86 netL86 6.828546707827616e-10
Rbbr86 netL86 0 -973287.030801482
Cbr86 netL86 0 1.1176275555033197e-21

* Branch 87
Rabr87 node_4 netRa87 6570168.227740637
Lbr87 netRa87 netL87 -1.205911117751876e-09
Rbbr87 netL87 0 -6899841.1271690875
Cbr87 netL87 0 -2.659998972602904e-23

* Branch 88
Rabr88 node_4 netRa88 -133015.9326049837
Lbr88 netRa88 netL88 1.018347964696193e-10
Rbbr88 netL88 0 345889.8895621987
Cbr88 netL88 0 2.2128146033696926e-21

* Branch 89
Rabr89 node_4 netRa89 152787.20944060612
Lbr89 netRa89 netL89 3.2693830158471234e-10
Rbbr89 netL89 0 -1525432.5343062533
Cbr89 netL89 0 1.403760793222098e-21

* Branch 90
Rabr90 node_4 netRa90 1069543.132914817
Lbr90 netRa90 netL90 4.40700820637107e-10
Rbbr90 netL90 0 -1389994.9034881743
Cbr90 netL90 0 2.96477677860615e-22

* Branch 91
Rabr91 node_4 netRa91 5740712.676460097
Lbr91 netRa91 netL91 8.753896674550123e-10
Rbbr91 netL91 0 -5957461.607748775
Cbr91 netL91 0 2.5597484996086102e-23

* Branch 92
Rabr92 node_4 netRa92 79323.41613321082
Lbr92 netRa92 netL92 1.7373640208267527e-10
Rbbr92 netL92 0 -769701.2140569738
Cbr92 netL92 0 2.8479349699359583e-21

* Branch 93
Rabr93 node_4 netRa93 82926.99671670959
Lbr93 netRa93 netL93 2.721827267424084e-10
Rbbr93 netL93 0 -1928302.3432588999
Cbr93 netL93 0 1.7046765436615622e-21

* Branch 94
Rabr94 node_4 netRa94 -55239.59573822552
Lbr94 netRa94 netL94 2.266632191614137e-10
Rbbr94 netL94 0 2756013.445752492
Cbr94 netL94 0 1.485999045012249e-21

* Branch 95
Rabr95 node_4 netRa95 168672.23673986315
Lbr95 netRa95 netL95 2.0263321243555032e-10
Rbbr95 netL95 0 -709394.7415478651
Cbr95 netL95 0 1.6947360525306385e-21

* Branch 96
Rabr96 node_4 netRa96 371584.82745167107
Lbr96 netRa96 netL96 4.1864059615063923e-10
Rbbr96 netL96 0 -1576533.4044426735
Cbr96 netL96 0 7.1516966356384085e-22

* Branch 97
Rabr97 node_4 netRa97 47065.12459628067
Lbr97 netRa97 netL97 1.225236423188521e-10
Rbbr97 netL97 0 -773713.5225327958
Cbr97 netL97 0 3.3712588999630465e-21

* Branch 98
Rabr98 node_4 netRa98 -38041.94638188566
Lbr98 netRa98 netL98 5.057286874246764e-11
Rbbr98 netL98 0 254762.65863486708
Cbr98 netL98 0 5.21240848009857e-21

* Branch 99
Rabr99 node_4 netRa99 -29826.611966359742
Lbr99 netRa99 netL99 -2.9943348908601825e-11
Rbbr99 netL99 0 136921.10165275115
Cbr99 netL99 0 -7.414243047004415e-21

.ends


.end
