* netlist generated with vector fitting poles and residues

.subckt total_network node_1 node_2 node_3 node_4 
X_11 node_1 0 yp11
X_12 node_1 node_2 yp12
X_13 node_1 node_3 yp13
X_14 node_1 node_4 yp14
X_22 node_2 0 yp22
X_23 node_2 node_3 yp23
X_24 node_2 node_4 yp24
X_33 node_3 0 yp33
X_34 node_3 node_4 yp34
X_44 node_4 0 yp44
.ends


* Y'11
.subckt yp11 node_1 0
* Branch 0
Rabr0 node_1 netRa0 -7.958350840997372
Lbr0 netRa0 netL0 -1.1830781945885065e-14
Rbbr0 netL0 0 18.480686487332108
Cbr0 netL0 0 -1.0265924759775643e-16

* Branch 1
Rabr1 node_1 netRa1 -9.547000796032664
Lbr1 netRa1 netL1 -2.0462890393332578e-14
Rbbr1 netL1 0 38.30791978553425
Cbr1 netL1 0 -7.848064479213709e-17

* Branch 2
Rabr2 node_1 netRa2 29.660751149527073
Lbr2 netRa2 netL2 5.567332836614375e-14
Rbbr2 netL2 0 -92.16072618896987
Cbr2 netL2 0 2.6111049786766096e-17

* Branch 3
Rabr3 node_1 netRa3 -1.4955344832506823
Lbr3 netRa3 netL3 1.1845833478325627e-14
Rbbr3 netL3 0 26.67574932531169
Cbr3 netL3 0 1.6825591969860572e-16

* Branch 4
Rabr4 node_1 netRa4 18.7390095532832
Lbr4 netRa4 netL4 -2.200650240562563e-14
Rbbr4 netL4 0 -30.326081487126736
Cbr4 netL4 0 -3.6317273357725894e-17

* Branch 5
Rabr5 node_1 netRa5 16.26710689939542
Lbr5 netRa5 netL5 -2.7095295741490392e-14
Rbbr5 netL5 0 -37.69947520250933
Cbr5 netL5 0 -4.108380802728898e-17

* Branch 6
Rabr6 node_1 netRa6 118.351027863159
Lbr6 netRa6 netL6 -1.795266720448153e-13
Rbbr6 netL6 0 -232.65152957858172
Cbr6 netL6 0 -6.138460184620919e-18

* Branch 7
Rabr7 node_1 netRa7 -211472.7658854312
Lbr7 netRa7 netL7 -2.4237976027954514e-11
Rbbr7 netL7 0 212602.65711563829
Cbr7 netL7 0 -5.409109052142843e-22

* Branch 8
Rabr8 node_1 netRa8 53.53394572136277
Lbr8 netRa8 netL8 9.726560890464266e-14
Rbbr8 netL8 0 -154.7650925924621
Cbr8 netL8 0 1.2328355414907465e-17

* Branch 9
Rabr9 node_1 netRa9 2.7920478938638644
Lbr9 netRa9 netL9 -1.6387184921058104e-14
Rbbr9 netL9 0 -106.86558578614252
Cbr9 netL9 0 -4.7837870456957386e-17

* Branch 10
Rabr10 node_1 netRa10 -23.697521161904085
Lbr10 netRa10 netL10 6.13214538537524e-14
Rbbr10 netL10 0 423.38247836024397
Cbr10 netL10 0 5.744708138415952e-18

* Branch 11
Rabr11 node_1 netRa11 801.4739331763558
Lbr11 netRa11 netL11 -1.2707384197811613e-13
Rbbr11 netL11 0 -855.1948026999648
Cbr11 netL11 0 -1.8470991602844678e-19

* Branch 12
Rabr12 node_1 netRa12 -96.35893016869896
Lbr12 netRa12 netL12 1.9113732202650903e-13
Rbbr12 netL12 0 1064.4948155405039
Cbr12 netL12 0 1.7883153061199e-18

* Branch 13
Rabr13 node_1 netRa13 1706.4623176470718
Lbr13 netRa13 netL13 -1.179203100120588e-12
Rbbr13 netL13 0 -4095.968201148439
Cbr13 netL13 0 -1.663440388592695e-19

* Branch 14
Rabr14 node_1 netRa14 259.7431774345058
Lbr14 netRa14 netL14 -2.8322048401396036e-13
Rbbr14 netL14 0 -1074.3433558744946
Cbr14 netL14 0 -9.930693507077896e-19

* Branch 15
Rabr15 node_1 netRa15 2949.4321621005806
Lbr15 netRa15 netL15 2.279866236610326e-13
Rbbr15 netL15 0 -2971.271375867113
Cbr15 netL15 0 2.6055811678849677e-20

* Branch 16
Rabr16 node_1 netRa16 -45.312884749438815
Lbr16 netRa16 netL16 3.470146174361002e-14
Rbbr16 netL16 0 78.01680187020952
Cbr16 netL16 0 9.672540523614614e-18

* Branch 17
Rabr17 node_1 netRa17 24567.286888855524
Lbr17 netRa17 netL17 -1.5300912474542416e-11
Rbbr17 netL17 0 -47686.21400123367
Cbr17 netL17 0 -1.2916085681504447e-20

* Branch 18
Rabr18 node_1 netRa18 -80774.3552526048
Lbr18 netRa18 netL18 2.6788081188723272e-11
Rbbr18 netL18 0 111818.25233886958
Cbr18 netL18 0 2.9483398189280454e-21

* Branch 19
Rabr19 node_1 netRa19 -325.9557709978776
Lbr19 netRa19 netL19 -8.126458811124661e-14
Rbbr19 netL19 0 351.1491608773507
Cbr19 netL19 0 -7.130471725271953e-19

* Branch 20
Rabr20 node_1 netRa20 480.64291026911445
Lbr20 netRa20 netL20 3.492356673556951e-12
Rbbr20 netL20 0 -40510.534825760464
Cbr20 netL20 0 2.0496328875553726e-19

* Branch 21
Rabr21 node_1 netRa21 -119356.81532768498
Lbr21 netRa21 netL21 -9.921723475439083e-11
Rbbr21 netL21 0 192164.12290057822
Cbr21 netL21 0 -4.387181530011197e-21

* Branch 22
Rabr22 node_1 netRa22 22.66063811433702
Lbr22 netRa22 netL22 1.2800745816290323e-13
Rbbr22 netL22 0 -2388.7981548310668
Cbr22 netL22 0 2.5931179638072768e-18

* Branch 23
Rabr23 node_1 netRa23 -522.7808412739612
Lbr23 netRa23 netL23 -1.0685853050506917e-11
Rbbr23 netL23 0 233057.79280663808
Cbr23 netL23 0 -1.2578491239012903e-19

* Branch 24
Rabr24 node_1 netRa24 -11542.39987717671
Lbr24 netRa24 netL24 -1.620215336645429e-11
Rbbr24 netL24 0 66066.87876703734
Cbr24 netL24 0 -2.167305515129852e-20

* Branch 25
Rabr25 node_1 netRa25 24352.563707480364
Lbr25 netRa25 netL25 3.3369418292597e-11
Rbbr25 netL25 0 -174653.8346666256
Cbr25 netL25 0 7.99497656555551e-21

* Branch 26
Rabr26 node_1 netRa26 8802.165802264693
Lbr26 netRa26 netL26 1.1177864681503005e-12
Rbbr26 netL26 0 -9227.736902082155
Cbr26 netL26 0 1.378529683808992e-20

* Branch 27
Rabr27 node_1 netRa27 1266.933609467216
Lbr27 netRa27 netL27 -2.169042991967436e-12
Rbbr27 netL27 0 -5548.817044852457
Cbr27 netL27 0 -3.0163691854265153e-19

* Branch 28
Rabr28 node_1 netRa28 -965931.7074550565
Lbr28 netRa28 netL28 -1.2743767681824732e-10
Rbbr28 netL28 0 984169.8604684459
Cbr28 netL28 0 -1.3428799065002862e-22

* Branch 29
Rabr29 node_1 netRa29 -867.5449481435481
Lbr29 netRa29 netL29 9.30945287218803e-13
Rbbr29 netL29 0 2121.8367455738107
Cbr29 netL29 0 4.989815136390193e-19

* Branch 30
Rabr30 node_1 netRa30 184920.0871586301
Lbr30 netRa30 netL30 3.386358381326502e-11
Rbbr30 netL30 0 -187799.4202405553
Cbr30 netL30 0 9.773586415705232e-22

* Branch 31
Rabr31 node_1 netRa31 6485.067840816036
Lbr31 netRa31 netL31 -7.342240867588766e-12
Rbbr31 netL31 0 -27466.59258282131
Cbr31 netL31 0 -4.064707072771984e-20

* Branch 32
Rabr32 node_1 netRa32 -9023.55938032158
Lbr32 netRa32 netL32 -3.466203537210907e-11
Rbbr32 netL32 0 134820.1029308933
Cbr32 netL32 0 -2.9814707598323885e-20

* Branch 33
Rabr33 node_1 netRa33 -56236.363418616565
Lbr33 netRa33 netL33 -9.358813296005255e-11
Rbbr33 netL33 0 188899.17516569103
Cbr33 netL33 0 -8.981530942163712e-21

* Branch 34
Rabr34 node_1 netRa34 -19574.37043569401
Lbr34 netRa34 netL34 -1.710378744167395e-11
Rbbr34 netL34 0 35520.22417189599
Cbr34 netL34 0 -2.4843291900477445e-20

* Branch 35
Rabr35 node_1 netRa35 -63.10540501890019
Lbr35 netRa35 netL35 6.097017862347596e-14
Rbbr35 netL35 0 170.063716556393
Cbr35 netL35 0 5.623816759996663e-18

* Branch 36
Rabr36 node_1 netRa36 -18313168.461724065
Lbr36 netRa36 netL36 3.0399812102895766e-10
Rbbr36 netL36 0 18324686.238920897
Cbr36 netL36 0 9.057320605546641e-25

* Branch 37
Rabr37 node_1 netRa37 -402781.8435554207
Lbr37 netRa37 netL37 -1.5577032708558573e-10
Rbbr37 netL37 0 579456.0193996066
Cbr37 netL37 0 -6.69875550564155e-22

* Branch 38
Rabr38 node_1 netRa38 70.23956584178106
Lbr38 netRa38 netL38 -5.0214956362109344e-14
Rbbr38 netL38 0 -135.91307414717426
Cbr38 netL38 0 -5.224622041410371e-18

* Branch 39
Rabr39 node_1 netRa39 2946.348584279787
Lbr39 netRa39 netL39 1.5041603351704735e-12
Rbbr39 netL39 0 -3357.6934994853727
Cbr39 netL39 0 1.5276854008103075e-19

* Branch 40
Rabr40 node_1 netRa40 -7277.389187703382
Lbr40 netRa40 netL40 -4.848264735150266e-11
Rbbr40 netL40 0 1096400.4249807002
Cbr40 netL40 0 -6.459998362369965e-21

* Branch 41
Rabr41 node_1 netRa41 372.19807067377326
Lbr41 netRa41 netL41 -1.0632512638782372e-12
Rbbr41 netL41 0 -1904.9175349040172
Cbr41 netL41 0 -1.4624664707807206e-18

* Branch 42
Rabr42 node_1 netRa42 55868.84032372777
Lbr42 netRa42 netL42 -1.9172554512143216e-11
Rbbr42 netL42 0 -60479.60688540641
Cbr42 netL42 0 -5.658690709807397e-21

* Branch 43
Rabr43 node_1 netRa43 -4099.412375553267
Lbr43 netRa43 netL43 -7.171476063064179e-12
Rbbr43 netL43 0 13176.880451319255
Cbr43 netL43 0 -1.3461762392512071e-19

* Branch 44
Rabr44 node_1 netRa44 -532.6206133362379
Lbr44 netRa44 netL44 -3.1944166257039894e-12
Rbbr44 netL44 0 14045.098496984232
Cbr44 netL44 0 -4.479967563917894e-19

* Branch 45
Rabr45 node_1 netRa45 -5007700.648679972
Lbr45 netRa45 netL45 3.450047768533392e-10
Rbbr45 netL45 0 5021681.879079144
Cbr45 netL45 0 1.3712557522166272e-23

* Branch 46
Rabr46 node_1 netRa46 40687.53998263368
Lbr46 netRa46 netL46 4.2245261371337475e-11
Rbbr46 netL46 0 -162762.45328981182
Cbr46 netL46 0 6.427849564374902e-21

* Branch 47
Rabr47 node_1 netRa47 -86062.52616419266
Lbr47 netRa47 netL47 7.793133626522608e-12
Rbbr47 netL47 0 87075.17051366006
Cbr47 netL47 0 1.039249358783234e-21

* Branch 48
Rabr48 node_1 netRa48 10097.02235505686
Lbr48 netRa48 netL48 1.015768481767431e-11
Rbbr48 netL48 0 -36294.66939983797
Cbr48 netL48 0 2.7920082280677187e-20

* Branch 49
Rabr49 node_1 netRa49 4462.352313805508
Lbr49 netRa49 netL49 6.364274592902791e-12
Rbbr49 netL49 0 -19150.507528055805
Cbr49 netL49 0 7.524584058070262e-20

* Branch 50
Rabr50 node_1 netRa50 -30695.604290604755
Lbr50 netRa50 netL50 -3.752416820602612e-11
Rbbr50 netL50 0 74013.01003264282
Cbr50 netL50 0 -1.6659789025966233e-20

* Branch 51
Rabr51 node_1 netRa51 13099.239764874663
Lbr51 netRa51 netL51 -5.960564887445614e-11
Rbbr51 netL51 0 -220717.83603467504
Cbr51 netL51 0 -2.000127175124512e-20

* Branch 52
Rabr52 node_1 netRa52 -9563.793101048333
Lbr52 netRa52 netL52 -2.289255034772883e-11
Rbbr52 netL52 0 201496.89317556572
Cbr52 netL52 0 -1.207344501113908e-20

* Branch 53
Rabr53 node_1 netRa53 -26208.68330530019
Lbr53 netRa53 netL53 5.75145091014699e-12
Rbbr53 netL53 0 29028.90010589279
Cbr53 netL53 0 7.549675380200931e-21

* Branch 54
Rabr54 node_1 netRa54 -519.7468153625402
Lbr54 netRa54 netL54 9.13600049629304e-13
Rbbr54 netL54 0 4006.1047757972715
Cbr54 netL54 0 4.342717428655622e-19

* Branch 55
Rabr55 node_1 netRa55 104054.50185107134
Lbr55 netRa55 netL55 -1.5169209193757413e-11
Rbbr55 netL55 0 -105518.15545719078
Cbr55 netL55 0 -1.3804473541035114e-21

* Branch 56
Rabr56 node_1 netRa56 1025453.4144835678
Lbr56 netRa56 netL56 -1.5839012941502477e-10
Rbbr56 netL56 0 -1040851.3121584095
Cbr56 netL56 0 -1.4827727518435457e-22

* Branch 57
Rabr57 node_1 netRa57 249125.43563050422
Lbr57 netRa57 netL57 -1.3432643065755519e-11
Rbbr57 netL57 0 -250183.91590869977
Cbr57 netL57 0 -2.1545893297734194e-22

* Branch 58
Rabr58 node_1 netRa58 -4358.08111996593
Lbr58 netRa58 netL58 -1.8701891434013303e-12
Rbbr58 netL58 0 5779.88462707153
Cbr58 netL58 0 -7.438865226864517e-20

* Branch 59
Rabr59 node_1 netRa59 -46186.56991642629
Lbr59 netRa59 netL59 -8.050686317273029e-11
Rbbr59 netL59 0 161020.6423297105
Cbr59 netL59 0 -1.090913563812569e-20

* Branch 60
Rabr60 node_1 netRa60 508.49329604688234
Lbr60 netRa60 netL60 1.2209240634185161e-12
Rbbr60 netL60 0 -5767.151314452565
Cbr60 netL60 0 4.2078745061771866e-19

* Branch 61
Rabr61 node_1 netRa61 19498.578395087752
Lbr61 netRa61 netL61 -9.0122006959613e-12
Rbbr61 netL61 0 -26477.410069682723
Cbr61 netL61 0 -1.7424406270138235e-20

* Branch 62
Rabr62 node_1 netRa62 5080.976830569915
Lbr62 netRa62 netL62 -3.161961007087831e-12
Rbbr62 netL62 0 -8045.406896197097
Cbr62 netL62 0 -7.717133338717635e-20

* Branch 63
Rabr63 node_1 netRa63 -139176.82731994192
Lbr63 netRa63 netL63 8.545179405344329e-11
Rbbr63 netL63 0 192548.7900552267
Cbr63 netL63 0 3.181439957556378e-21

* Branch 64
Rabr64 node_1 netRa64 172969.50012324023
Lbr64 netRa64 netL64 -2.7357300399175316e-11
Rbbr64 netL64 0 -179701.63167516343
Cbr64 netL64 0 -8.796410105646842e-22

* Branch 65
Rabr65 node_1 netRa65 47047.2533034151
Lbr65 netRa65 netL65 1.9969677071010287e-11
Rbbr65 netL65 0 -73259.24322504157
Cbr65 netL65 0 5.801787107348278e-21

* Branch 66
Rabr66 node_1 netRa66 7633.942056390867
Lbr66 netRa66 netL66 -8.309764271372639e-12
Rbbr66 netL66 0 -26015.084235700273
Cbr66 netL66 0 -4.1698014511422774e-20

* Branch 67
Rabr67 node_1 netRa67 11915.921797703313
Lbr67 netRa67 netL67 1.5900372056291107e-11
Rbbr67 netL67 0 -76954.82581150424
Cbr67 netL67 0 1.7406804588447172e-20

* Branch 68
Rabr68 node_1 netRa68 -554.2008165478196
Lbr68 netRa68 netL68 4.120456124380249e-13
Rbbr68 netL68 0 1119.2211553430784
Cbr68 netL68 0 6.6311036466600515e-19

* Branch 69
Rabr69 node_1 netRa69 -808808.5539048009
Lbr69 netRa69 netL69 1.3056062943175e-10
Rbbr69 netL69 0 829806.4526740481
Cbr69 netL69 0 1.9447919685321775e-22

* Branch 70
Rabr70 node_1 netRa70 -315126.6832452109
Lbr70 netRa70 netL70 7.298839771758624e-11
Rbbr70 netL70 0 331333.47932486737
Cbr70 netL70 0 6.988002301398163e-22

* Branch 71
Rabr71 node_1 netRa71 -3355308.6205214257
Lbr71 netRa71 netL71 3.2880261220575903e-10
Rbbr71 netL71 0 3432178.579370603
Cbr71 netL71 0 2.8547744199075606e-23

* Branch 72
Rabr72 node_1 netRa72 194044.4712411718
Lbr72 netRa72 netL72 2.336392419902636e-11
Rbbr72 netL72 0 -199720.41047103461
Cbr72 netL72 0 6.029679210039228e-22

* Branch 73
Rabr73 node_1 netRa73 1856575.3398323418
Lbr73 netRa73 netL73 6.357399568792132e-11
Rbbr73 netL73 0 -1860186.9722133758
Cbr73 netL73 0 1.840892979364147e-23

* Branch 74
Rabr74 node_1 netRa74 -30665.497195858687
Lbr74 netRa74 netL74 -2.435111001040111e-11
Rbbr74 netL74 0 71491.86530429452
Cbr74 netL74 0 -1.1117188696794369e-20

* Branch 75
Rabr75 node_1 netRa75 -709718.713543705
Lbr75 netRa75 netL75 2.340395931782244e-10
Rbbr75 netL75 0 927887.1626070355
Cbr75 netL75 0 3.5526387832114097e-22

* Branch 76
Rabr76 node_1 netRa76 -249496.22887796094
Lbr76 netRa76 netL76 2.944092887617253e-11
Rbbr76 netL76 0 256268.4719458382
Cbr76 netL76 0 4.60402625340158e-22

* Branch 77
Rabr77 node_1 netRa77 755566.7155096444
Lbr77 netRa77 netL77 1.0912483350169404e-10
Rbbr77 netL77 0 -805087.2656818511
Cbr77 netL77 0 1.7941544133160316e-22

* Branch 78
Rabr78 node_1 netRa78 -506616.3096089396
Lbr78 netRa78 netL78 1.0950345017513824e-10
Rbbr78 netL78 0 584671.9284293827
Cbr78 netL78 0 3.6965630231137423e-22

* Branch 79
Rabr79 node_1 netRa79 -1727996.5833456728
Lbr79 netRa79 netL79 -1.7344144683356414e-10
Rbbr79 netL79 0 1764092.3064221907
Cbr79 netL79 0 -5.689751799954739e-23

* Branch 80
Rabr80 node_1 netRa80 -1456222.342318971
Lbr80 netRa80 netL80 1.1000267526506245e-10
Rbbr80 netL80 0 1464382.704995948
Cbr80 netL80 0 5.1583050944169144e-23

* Branch 81
Rabr81 node_1 netRa81 -650708.7476811704
Lbr81 netRa81 netL81 -3.156635548940639e-10
Rbbr81 netL81 0 1030727.8359938057
Cbr81 netL81 0 -4.70754767161785e-22

* Branch 82
Rabr82 node_1 netRa82 -5703622.999366024
Lbr82 netRa82 netL82 4.2392590605378675e-10
Rbbr82 netL82 0 5809159.837460132
Cbr82 netL82 0 1.2794090185840703e-23

* Branch 83
Rabr83 node_1 netRa83 -62389.895902451266
Lbr83 netRa83 netL83 1.046715822826544e-11
Rbbr83 netL83 0 65751.53200429189
Cbr83 netL83 0 2.551125792220248e-21

* Branch 84
Rabr84 node_1 netRa84 9161292.419616172
Lbr84 netRa84 netL84 2.922225815546937e-10
Rbbr84 netL84 0 -9176513.963197125
Cbr84 netL84 0 3.476114611214238e-24

* Branch 85
Rabr85 node_1 netRa85 155138.13106895424
Lbr85 netRa85 netL85 5.248906964254463e-11
Rbbr85 netL85 0 -175380.92700151843
Cbr85 netL85 0 1.9298636688386054e-21

* Branch 86
Rabr86 node_1 netRa86 28125.445668318494
Lbr86 netRa86 netL86 3.3357021622096134e-11
Rbbr86 netL86 0 -74176.1242031911
Cbr86 netL86 0 1.601104349780412e-20

* Branch 87
Rabr87 node_1 netRa87 16290.408297728574
Lbr87 netRa87 netL87 -5.044772708093345e-12
Rbbr87 netL87 0 -18623.051761304392
Cbr87 netL87 0 -1.6622633042718454e-20

* Branch 88
Rabr88 node_1 netRa88 -96.28949684316906
Lbr88 netRa88 netL88 7.497844843471296e-13
Rbbr88 netL88 0 8410.131689461441
Cbr88 netL88 0 9.132891805571583e-19

* Branch 89
Rabr89 node_1 netRa89 -4316.729613995331
Lbr89 netRa89 netL89 1.5678422028081604e-12
Rbbr89 netL89 0 5385.148490622405
Cbr89 netL89 0 6.739997159923441e-20

* Branch 90
Rabr90 node_1 netRa90 -3276.1387568621503
Lbr90 netRa90 netL90 -1.2233334877319817e-12
Rbbr90 netL90 0 4291.4048286437355
Cbr90 netL90 0 -8.710967080566212e-20

* Branch 91
Rabr91 node_1 netRa91 631.1835216203341
Lbr91 netRa91 netL91 6.742937609841051e-12
Rbbr91 netL91 0 -49975.53728693269
Cbr91 netL91 0 2.239408392445894e-19

* Branch 92
Rabr92 node_1 netRa92 -787682.5280986882
Lbr92 netRa92 netL92 -6.809525529519165e-11
Rbbr92 netL92 0 808197.5539229708
Cbr92 netL92 0 -1.07007902326874e-22

* Branch 93
Rabr93 node_1 netRa93 4288.200369765463
Lbr93 netRa93 netL93 -1.0537837750345305e-12
Rbbr93 netL93 0 -4857.760597839043
Cbr93 netL93 0 -5.051415287384464e-20

* Branch 94
Rabr94 node_1 netRa94 27967.486972860548
Lbr94 netRa94 netL94 2.5112759746778777e-11
Rbbr94 netL94 0 -58381.82277856726
Cbr94 netL94 0 1.5490645166364416e-20

* Branch 95
Rabr95 node_1 netRa95 -159.33136879903728
Lbr95 netRa95 netL95 -1.2477939494903299e-13
Rbbr95 netL95 0 455.08006554181304
Cbr95 netL95 0 -1.7439219914848887e-18

* Branch 96
Rabr96 node_1 netRa96 -390.76686856922055
Lbr96 netRa96 netL96 -9.35253653963157e-14
Rbbr96 netL96 0 451.1154466894343
Cbr96 netL96 0 -5.339963896430529e-19

* Branch 97
Rabr97 node_1 netRa97 -54.04649690938559
Lbr97 netRa97 netL97 -4.529626733916044e-14
Rbbr97 netL97 0 74.97220531363128
Cbr97 netL97 0 -1.1501268143780912e-17

* Branch 98
Rabr98 node_1 netRa98 10.597947989483272
Lbr98 netRa98 netL98 2.397205493491878e-14
Rbbr98 netL98 0 -84.55077472290148
Cbr98 netL98 0 2.912107291109014e-17

* Branch 99
Rabr99 node_1 netRa99 1.8132336167536371
Lbr99 netRa99 netL99 7.800492658965758e-15
Rbbr99 netL99 0 -27.9662549737644
Cbr99 netL99 0 2.603765122739878e-16

.ends


* Y'12
.subckt yp12 node_1 node_2
* Branch 0
Rabr0 node_1 netRa0 544.2747355865685
Lbr0 netRa0 netL0 -8.701265092418646e-14
Rbbr0 netL0 node_2 -554.2316865416359
Cbr0 netL0 node_2 -2.8370565128549e-19

* Branch 1
Rabr1 node_1 netRa1 247.71725758326335
Lbr1 netRa1 netL1 5.236409739129229e-14
Rbbr1 netL1 node_2 -255.9319051541789
Cbr1 netL1 node_2 8.435678798840945e-19

* Branch 2
Rabr2 node_1 netRa2 27.435764484710173
Lbr2 netRa2 netL2 1.835693723445052e-14
Rbbr2 netL2 node_2 -36.99380749582263
Cbr2 netL2 node_2 1.930118464256721e-17

* Branch 3
Rabr3 node_1 netRa3 2.8640901639134446
Lbr3 netRa3 netL3 7.358294704315974e-15
Rbbr3 netL3 node_2 -20.391915081481173
Cbr3 netL3 node_2 1.5937878924985526e-16

* Branch 4
Rabr4 node_1 netRa4 4.84947216805926
Lbr4 netRa4 netL4 1.6763656910793183e-14
Rbbr4 netL4 node_2 -44.24729781266852
Cbr4 netL4 node_2 1.0223203076193158e-16

* Branch 5
Rabr5 node_1 netRa5 -118.67460001784872
Lbr5 netRa5 netL5 2.1863738868954913e-13
Rbbr5 netL5 node_2 271.90932966994006
Cbr5 netL5 node_2 6.1970912200346486e-18

* Branch 6
Rabr6 node_1 netRa6 31.995405253969842
Lbr6 netRa6 netL6 -3.687504326394836e-14
Rbbr6 netL6 node_2 -149.4145023416816
Cbr6 netL6 node_2 -7.304534158486406e-18

* Branch 7
Rabr7 node_1 netRa7 -0.35912977563210446
Lbr7 netRa7 netL7 -3.881131557006913e-15
Rbbr7 netL7 node_2 50.745730339489754
Cbr7 netL7 node_2 -3.3540272680647357e-16

* Branch 8
Rabr8 node_1 netRa8 72.46483669699478
Lbr8 netRa8 netL8 -3.053544013606199e-14
Rbbr8 netL8 node_2 -106.61018310176883
Cbr8 netL8 node_2 -3.899890325573887e-18

* Branch 9
Rabr9 node_1 netRa9 1448.4212660393985
Lbr9 netRa9 netL9 -2.7145359033868748e-12
Rbbr9 netL9 node_2 -17750.840345173143
Cbr9 netL9 node_2 -9.971703929438388e-20

* Branch 10
Rabr10 node_1 netRa10 15.346845120798536
Lbr10 netRa10 netL10 1.4931289736919934e-14
Rbbr10 netL10 node_2 -48.520976403560304
Cbr10 netL10 node_2 2.0631243840020292e-17

* Branch 11
Rabr11 node_1 netRa11 119.02190648147024
Lbr11 netRa11 netL11 4.4134180240305676e-14
Rbbr11 netL11 node_2 -158.99156234464172
Cbr11 netL11 node_2 2.3559052421532287e-18

* Branch 12
Rabr12 node_1 netRa12 -5692.925507374005
Lbr12 netRa12 netL12 5.5368721311029265e-12
Rbbr12 netL12 node_2 22945.498547951847
Cbr12 netL12 node_2 4.1331816254992024e-20

* Branch 13
Rabr13 node_1 netRa13 4.733234144530969
Lbr13 netRa13 netL13 8.03896500664284e-15
Rbbr13 netL13 node_2 -35.05527411997518
Cbr13 netL13 node_2 5.0675349755716905e-17

* Branch 14
Rabr14 node_1 netRa14 15.139095974418654
Lbr14 netRa14 netL14 -1.8131928636766412e-14
Rbbr14 netL14 node_2 -69.14400327011134
Cbr14 netL14 node_2 -1.6812286022896532e-17

* Branch 15
Rabr15 node_1 netRa15 9.440973437798275
Lbr15 netRa15 netL15 -5.0313634660852596e-14
Rbbr15 netL15 node_2 -720.6231640954699
Cbr15 netL15 node_2 -6.53540432357486e-18

* Branch 16
Rabr16 node_1 netRa16 -87.04326910357553
Lbr16 netRa16 netL16 4.863339470880984e-14
Rbbr16 netL16 node_2 167.8634037787314
Cbr16 netL16 node_2 3.283643695909525e-18

* Branch 17
Rabr17 node_1 netRa17 690.4219307316184
Lbr17 netRa17 netL17 1.4769526633854164e-13
Rbbr17 netL17 node_2 -785.9209495383784
Cbr17 netL17 node_2 2.7360842402155546e-19

* Branch 18
Rabr18 node_1 netRa18 -14.141870020079129
Lbr18 netRa18 netL18 2.0026598618067633e-14
Rbbr18 netL18 node_2 64.62649100224819
Cbr18 netL18 node_2 2.1191528991564676e-17

* Branch 19
Rabr19 node_1 netRa19 23.00697087833893
Lbr19 netRa19 netL19 1.5992440344197206e-14
Rbbr19 netL19 node_2 -51.63328261952103
Cbr19 netL19 node_2 1.3689402979825092e-17

* Branch 20
Rabr20 node_1 netRa20 482.6218718940859
Lbr20 netRa20 netL20 7.328057198085248e-14
Rbbr20 netL20 node_2 -507.86743994242295
Cbr20 netL20 node_2 3.0003946921387533e-19

* Branch 21
Rabr21 node_1 netRa21 131.54212710227353
Lbr21 netRa21 netL21 -6.640341669689147e-14
Rbbr21 netL21 node_2 -168.28330390231127
Cbr21 netL21 node_2 -2.965963932032328e-18

* Branch 22
Rabr22 node_1 netRa22 -13.9209690201864
Lbr22 netRa22 netL22 -4.236581471368121e-14
Rbbr22 netL22 node_2 138.8544550158743
Cbr22 netL22 node_2 -2.352439755950887e-17

* Branch 23
Rabr23 node_1 netRa23 38.9257407566365
Lbr23 netRa23 netL23 2.949077447346402e-14
Rbbr23 netL23 node_2 -88.21748245486634
Cbr23 netL23 node_2 8.7337600927417e-18

* Branch 24
Rabr24 node_1 netRa24 -15.22384403162685
Lbr24 netRa24 netL24 1.610260144821364e-14
Rbbr24 netL24 node_2 39.59318713661025
Cbr24 netL24 node_2 2.611640098470667e-17

* Branch 25
Rabr25 node_1 netRa25 37.02959700159177
Lbr25 netRa25 netL25 5.1657080287580656e-14
Rbbr25 netL25 node_2 -263.15598248599196
Cbr25 netL25 node_2 5.465433991529576e-18

* Branch 26
Rabr26 node_1 netRa26 -15.095349362505068
Lbr26 netRa26 netL26 1.1106097876672225e-14
Rbbr26 netL26 node_2 26.566811265433554
Cbr26 netL26 node_2 2.7262529255043945e-17

* Branch 27
Rabr27 node_1 netRa27 -8.807322293046004
Lbr27 netRa27 netL27 -2.6592483334879514e-14
Rbbr27 netL27 node_2 79.438547796933
Cbr27 netL27 node_2 -4.0623513179189805e-17

* Branch 28
Rabr28 node_1 netRa28 -442.2346616084297
Lbr28 netRa28 netL28 4.444038435449675e-13
Rbbr28 netL28 node_2 1801.3268667525606
Cbr28 netL28 node_2 5.465552679018862e-19

* Branch 29
Rabr29 node_1 netRa29 -12.24895931951207
Lbr29 netRa29 netL29 1.8822807193570182e-14
Rbbr29 netL29 node_2 65.83546232211303
Cbr29 netL29 node_2 2.2625658931839048e-17

* Branch 30
Rabr30 node_1 netRa30 92.27996128844991
Lbr30 netRa30 netL30 -7.243979472683415e-14
Rbbr30 netL30 node_2 -152.39619867994486
Cbr30 netL30 node_2 -5.069466339861556e-18

* Branch 31
Rabr31 node_1 netRa31 496.7940070272497
Lbr31 netRa31 netL31 7.837904743562032e-14
Rbbr31 netL31 node_2 -511.0702672331564
Cbr31 netL31 node_2 3.097031670981125e-19

* Branch 32
Rabr32 node_1 netRa32 -2.2124162636849456
Lbr32 netRa32 netL32 2.1861635352274313e-14
Rbbr32 netL32 node_2 353.03644110957066
Cbr32 netL32 node_2 2.3314959456817258e-17

* Branch 33
Rabr33 node_1 netRa33 -1.8093467796113571
Lbr33 netRa33 netL33 2.5641471234862466e-14
Rbbr33 netL33 node_2 568.1722853642924
Cbr33 netL33 node_2 1.9518217932950883e-17

* Branch 34
Rabr34 node_1 netRa34 227.36906984113995
Lbr34 netRa34 netL34 -1.2340958091584487e-13
Rbbr34 netL34 node_2 -296.6725305942684
Cbr34 netL34 node_2 -1.810796595486539e-18

* Branch 35
Rabr35 node_1 netRa35 2.8779872501142187
Lbr35 netRa35 netL35 -6.294702145749612e-14
Rbbr35 netL35 node_2 -690.6186996745571
Cbr35 netL35 node_2 -2.2420238182740325e-17

* Branch 36
Rabr36 node_1 netRa36 -44.50841623446919
Lbr36 netRa36 netL36 -5.087312499486561e-14
Rbbr36 netL36 node_2 94.77790590001074
Cbr36 netL36 node_2 -1.2320239405986887e-17

* Branch 37
Rabr37 node_1 netRa37 -53.35359511878492
Lbr37 netRa37 netL37 1.54953759332125e-14
Rbbr37 netL37 node_2 59.58543467630422
Cbr37 netL37 node_2 4.84867181802339e-18

* Branch 38
Rabr38 node_1 netRa38 -43.66558810106286
Lbr38 netRa38 netL38 -6.822381077310312e-14
Rbbr38 netL38 node_2 139.33815661421852
Cbr38 netL38 node_2 -1.1531326816320797e-17

* Branch 39
Rabr39 node_1 netRa39 534.5133762568618
Lbr39 netRa39 netL39 -1.596107108259127e-13
Rbbr39 netL39 node_2 -650.7367975964903
Cbr39 netL39 node_2 -4.5648634184798925e-19

* Branch 40
Rabr40 node_1 netRa40 -42.56622850500029
Lbr40 netRa40 netL40 -7.715454563156544e-14
Rbbr40 netL40 node_2 176.88838354677623
Cbr40 netL40 node_2 -1.0577279879746422e-17

* Branch 41
Rabr41 node_1 netRa41 208.7057909027028
Lbr41 netRa41 netL41 -1.616885226551015e-13
Rbbr41 netL41 node_2 -555.0622620191373
Cbr41 netL41 node_2 -1.3776503486147657e-18

* Branch 42
Rabr42 node_1 netRa42 -31.139164724026408
Lbr42 netRa42 netL42 3.8380556724475155e-14
Rbbr42 netL42 node_2 114.6326259847662
Cbr42 netL42 node_2 1.0538878280551095e-17

* Branch 43
Rabr43 node_1 netRa43 972.0256125473829
Lbr43 netRa43 netL43 -2.6913584350762843e-13
Rbbr43 netL43 node_2 -1166.6322358957393
Cbr43 netL43 node_2 -2.362658096264292e-19

* Branch 44
Rabr44 node_1 netRa44 366.3054732537187
Lbr44 netRa44 netL44 1.3803720148578895e-13
Rbbr44 netL44 node_2 -490.2980999733956
Cbr44 netL44 node_2 7.732347183289479e-19

* Branch 45
Rabr45 node_1 netRa45 -514.4326453127089
Lbr45 netRa45 netL45 -1.440696841101754e-13
Rbbr45 netL45 node_2 546.4904729284866
Cbr45 netL45 node_2 -5.146809509421912e-19

* Branch 46
Rabr46 node_1 netRa46 -14.038084677035263
Lbr46 netRa46 netL46 2.969994852138887e-14
Rbbr46 netL46 node_2 121.33923098325607
Cbr46 netL46 node_2 1.689302592212043e-17

* Branch 47
Rabr47 node_1 netRa47 97.96690785388404
Lbr47 netRa47 netL47 -1.2944958506079387e-13
Rbbr47 netL47 node_2 -267.8302104717362
Cbr47 netL47 node_2 -4.8373343186819316e-18

* Branch 48
Rabr48 node_1 netRa48 -114.88291561682696
Lbr48 netRa48 netL48 -3.372505178620811e-14
Rbbr48 netL48 node_2 129.98069278807668
Cbr48 netL48 node_2 -2.2684570490744007e-18

* Branch 49
Rabr49 node_1 netRa49 45087.6230732605
Lbr49 netRa49 netL49 -1.2199041365867012e-12
Rbbr49 netL49 node_2 -45164.241405865025
Cbr49 netL49 node_2 -5.988264494028296e-22

* Branch 50
Rabr50 node_1 netRa50 -97.69175544799582
Lbr50 netRa50 netL50 3.762450671614743e-14
Rbbr50 netL50 node_2 127.9698559500849
Cbr50 netL50 node_2 2.992800159566525e-18

* Branch 51
Rabr51 node_1 netRa51 -6.963791194525757
Lbr51 netRa51 netL51 1.930913657562485e-14
Rbbr51 netL51 node_2 95.75105497876092
Cbr51 netL51 node_2 2.783594523941074e-17

* Branch 52
Rabr52 node_1 netRa52 -411.57225963736283
Lbr52 netRa52 netL52 -1.8142835088017093e-13
Rbbr52 netL52 node_2 631.4665216346903
Cbr52 netL52 node_2 -7.025082023905467e-19

* Branch 53
Rabr53 node_1 netRa53 45.30670086731523
Lbr53 netRa53 netL53 -1.5070751417628264e-14
Rbbr53 netL53 node_2 -51.20122897222568
Cbr53 netL53 node_2 -6.466447858948732e-18

* Branch 54
Rabr54 node_1 netRa54 139.7916946174484
Lbr54 netRa54 netL54 -9.918906737989136e-14
Rbbr54 netL54 node_2 -190.96116823956584
Cbr54 netL54 node_2 -3.680895145932324e-18

* Branch 55
Rabr55 node_1 netRa55 -14.790091218430142
Lbr55 netRa55 netL55 1.8212696032979103e-14
Rbbr55 netL55 node_2 49.99674781441448
Cbr55 netL55 node_2 2.424572573945413e-17

* Branch 56
Rabr56 node_1 netRa56 -58.47210057605751
Lbr56 netRa56 netL56 3.5538633155864563e-14
Rbbr56 netL56 node_2 94.8850951027309
Cbr56 netL56 node_2 6.359581319607705e-18

* Branch 57
Rabr57 node_1 netRa57 4.349254440937208
Lbr57 netRa57 netL57 3.773345325140597e-14
Rbbr57 netL57 node_2 -279.91471266071244
Cbr57 netL57 node_2 3.4230021954290616e-17

* Branch 58
Rabr58 node_1 netRa58 -453.5128007978976
Lbr58 netRa58 netL58 1.5963940583251923e-13
Rbbr58 netL58 node_2 558.9694594997593
Cbr58 netL58 node_2 6.273924477921659e-19

* Branch 59
Rabr59 node_1 netRa59 -54.33872883475126
Lbr59 netRa59 netL59 -1.4818936932999572e-13
Rbbr59 netL59 node_2 452.7872394437128
Cbr59 netL59 node_2 -6.200636903987392e-18

* Branch 60
Rabr60 node_1 netRa60 -38.15562318748906
Lbr60 netRa60 netL60 2.5672187311127887e-14
Rbbr60 netL60 node_2 64.9763765023042
Cbr60 netL60 node_2 1.0282345993578783e-17

* Branch 61
Rabr61 node_1 netRa61 -45.19300297565159
Lbr61 netRa61 netL61 3.849396961644289e-14
Rbbr61 netL61 node_2 99.26755094190341
Cbr61 netL61 node_2 8.506333822633481e-18

* Branch 62
Rabr62 node_1 netRa62 -65.68657997507462
Lbr62 netRa62 netL62 7.19671316651569e-14
Rbbr62 netL62 node_2 224.35976706681774
Cbr62 netL62 node_2 4.829734162715021e-18

* Branch 63
Rabr63 node_1 netRa63 -22.169052555559645
Lbr63 netRa63 netL63 3.068947256149049e-14
Rbbr63 netL63 node_2 90.4266921435529
Cbr63 netL63 node_2 1.509917025556904e-17

* Branch 64
Rabr64 node_1 netRa64 -422.5566653962434
Lbr64 netRa64 netL64 -5.111561844254497e-14
Rbbr64 netL64 node_2 431.01030671835116
Cbr64 netL64 node_2 -2.8099540405790323e-19

* Branch 65
Rabr65 node_1 netRa65 -4.7971922334978405
Lbr65 netRa65 netL65 -1.7373004487759917e-13
Rbbr65 netL65 node_2 9330.119055707828
Cbr65 netL65 node_2 -5.851161646431647e-18

* Branch 66
Rabr66 node_1 netRa66 53134.2403153723
Lbr66 netRa66 netL66 5.862988289326852e-12
Rbbr66 netL66 node_2 -53515.70792425156
Cbr66 netL66 node_2 2.063903663557443e-21

* Branch 67
Rabr67 node_1 netRa67 -258.26302077068414
Lbr67 netRa67 netL67 -1.7045923197017088e-13
Rbbr67 netL67 node_2 544.0509009029315
Cbr67 netL67 node_2 -1.2198567536654785e-18

* Branch 68
Rabr68 node_1 netRa68 427.3081960514305
Lbr68 netRa68 netL68 2.213674727998157e-12
Rbbr68 netL68 node_2 -39068.81494749189
Cbr68 netL68 node_2 1.3825118757765606e-19

* Branch 69
Rabr69 node_1 netRa69 -145.3933924238648
Lbr69 netRa69 netL69 9.32621049058489e-14
Rbbr69 netL69 node_2 268.603146649234
Cbr69 netL69 node_2 2.377116771568041e-18

* Branch 70
Rabr70 node_1 netRa70 -1528.3116542942662
Lbr70 netRa70 netL70 -1.2126910209475222e-12
Rbbr70 netL70 node_2 2179.8508260983936
Cbr70 netL70 node_2 -3.6608172591982257e-19

* Branch 71
Rabr71 node_1 netRa71 -92656.36760354678
Lbr71 netRa71 netL71 1.0130410548214225e-11
Rbbr71 netL71 node_2 96159.41415742939
Cbr71 netL71 node_2 1.136113204074426e-21

* Branch 72
Rabr72 node_1 netRa72 -203343.6014751716
Lbr72 netRa72 netL72 5.850147492158848e-12
Rbbr72 netL72 node_2 203796.98420529542
Cbr72 netL72 node_2 1.411418610954044e-22

* Branch 73
Rabr73 node_1 netRa73 2416.5642589940794
Lbr73 netRa73 netL73 1.959965373230914e-12
Rbbr73 netL73 node_2 -3393.9901193906185
Cbr73 netL73 node_2 2.402055631338068e-19

* Branch 74
Rabr74 node_1 netRa74 -469.1124781356382
Lbr74 netRa74 netL74 9.552773314732954e-13
Rbbr74 netL74 node_2 1703.528037155525
Cbr74 netL74 node_2 1.180939553764455e-18

* Branch 75
Rabr75 node_1 netRa75 -1.5385921835876912
Lbr75 netRa75 netL75 -9.617882700244224e-15
Rbbr75 netL75 node_2 79.08093878446708
Cbr75 netL75 node_2 -8.19969977550805e-17

* Branch 76
Rabr76 node_1 netRa76 25900.22094456982
Lbr76 netRa76 netL76 -1.4738409713846424e-12
Rbbr76 netL76 node_2 -26092.162185406458
Cbr76 netL76 node_2 -2.1802375108305806e-21

* Branch 77
Rabr77 node_1 netRa77 -70.98544334269937
Lbr77 netRa77 netL77 5.644071916102165e-14
Rbbr77 netL77 node_2 139.58261261801164
Cbr77 netL77 node_2 5.672962749998633e-18

* Branch 78
Rabr78 node_1 netRa78 910.9682538922194
Lbr78 netRa78 netL78 -6.644052335992094e-13
Rbbr78 netL78 node_2 -2566.1140744995173
Cbr78 netL78 node_2 -2.8316735714628184e-19

* Branch 79
Rabr79 node_1 netRa79 959.7457297025205
Lbr79 netRa79 netL79 -1.4508008335921085e-12
Rbbr79 netL79 node_2 -7214.767737692977
Cbr79 netL79 node_2 -2.0803745558897609e-19

* Branch 80
Rabr80 node_1 netRa80 1444.6697962035553
Lbr80 netRa80 netL80 -1.280361733621502e-12
Rbbr80 netL80 node_2 -2085.652955441977
Cbr80 netL80 node_2 -4.231745273099356e-19

* Branch 81
Rabr81 node_1 netRa81 455.1901173384819
Lbr81 netRa81 netL81 -1.1984801392310881e-12
Rbbr81 netL81 node_2 -9312.98133278145
Cbr81 netL81 node_2 -2.8003097350929896e-19

* Branch 82
Rabr82 node_1 netRa82 -9.790059455306382
Lbr82 netRa82 netL82 -1.6662944757386616e-14
Rbbr82 netL82 node_2 44.4450616055101
Cbr82 netL82 node_2 -3.8519495809116363e-17

* Branch 83
Rabr83 node_1 netRa83 -254745.90360837098
Lbr83 netRa83 netL83 8.065865749238182e-12
Rbbr83 netL83 node_2 255673.8451362954
Cbr83 netL83 node_2 1.2382741855758788e-22

* Branch 84
Rabr84 node_1 netRa84 -3.549281804542654
Lbr84 netRa84 netL84 -5.041241481125711e-15
Rbbr84 netL84 node_2 13.004141228898371
Cbr84 netL84 node_2 -1.0967804908378646e-16

* Branch 85
Rabr85 node_1 netRa85 -1.250764285674678
Lbr85 netRa85 netL85 -9.18684207267222e-15
Rbbr85 netL85 node_2 89.00310392648574
Cbr85 netL85 node_2 -8.424940382115585e-17

* Branch 86
Rabr86 node_1 netRa86 -0.4540117076704194
Lbr86 netRa86 netL86 -2.9698552674794314e-15
Rbbr86 netL86 node_2 26.144174642304876
Cbr86 netL86 node_2 -2.548445981571939e-16

* Branch 87
Rabr87 node_1 netRa87 -14.486622151354574
Lbr87 netRa87 netL87 1.2131263223092752e-14
Rbbr87 netL87 node_2 28.023518138226596
Cbr87 netL87 node_2 2.981551075257381e-17

* Branch 88
Rabr88 node_1 netRa88 9.748793670968926
Lbr88 netRa88 netL88 -2.4049511008003756e-14
Rbbr88 netL88 node_2 -80.04019890358077
Cbr88 netL88 node_2 -3.06294568663462e-17

* Branch 89
Rabr89 node_1 netRa89 -793.0139056566635
Lbr89 netRa89 netL89 -1.0670637071154602e-12
Rbbr89 netL89 node_2 1499.580276343299
Cbr89 netL89 node_2 -9.001583597983271e-19

* Branch 90
Rabr90 node_1 netRa90 -611.6264333082726
Lbr90 netRa90 netL90 -9.458175870514116e-13
Rbbr90 netL90 node_2 1358.5528354322942
Cbr90 netL90 node_2 -1.1422581529186415e-18

* Branch 91
Rabr91 node_1 netRa91 1855.4892695041149
Lbr91 netRa91 netL91 2.782908532981679e-12
Rbbr91 netL91 node_2 -15249.188944222751
Cbr91 netL91 node_2 9.867533289373226e-20

* Branch 92
Rabr92 node_1 netRa92 -302.83252225360803
Lbr92 netRa92 netL92 -1.2967617275103827e-12
Rbbr92 netL92 node_2 3355.724693190915
Cbr92 netL92 node_2 -1.2822178202957766e-18

* Branch 93
Rabr93 node_1 netRa93 -1189.299224869727
Lbr93 netRa93 netL93 -1.572266425975408e-12
Rbbr93 netL93 node_2 2287.7995043151577
Cbr93 netL93 node_2 -5.786468879646607e-19

* Branch 94
Rabr94 node_1 netRa94 -729.5340280505752
Lbr94 netRa94 netL94 -1.1680881367561593e-12
Rbbr94 netL94 node_2 1613.8110088228816
Cbr94 netL94 node_2 -9.934109628043754e-19

* Branch 95
Rabr95 node_1 netRa95 -387.7669603557341
Lbr95 netRa95 netL95 -4.834219697080103e-13
Rbbr95 netL95 node_2 657.1529756375719
Cbr95 netL95 node_2 -1.8984898715402984e-18

* Branch 96
Rabr96 node_1 netRa96 -505.3002776813186
Lbr96 netRa96 netL96 5.941425920853926e-13
Rbbr96 netL96 node_2 821.60556933573
Cbr96 netL96 node_2 1.426145061521741e-18

* Branch 97
Rabr97 node_1 netRa97 -945.4883315709437
Lbr97 netRa97 netL97 5.927916971535738e-13
Rbbr97 netL97 node_2 2213.830043993607
Cbr97 netL97 node_2 2.8182697552071885e-19

* Branch 98
Rabr98 node_1 netRa98 -22.902086838722234
Lbr98 netRa98 netL98 -2.3206810502790538e-14
Rbbr98 netL98 node_2 96.29988799997419
Cbr98 netL98 node_2 -1.0849461254883325e-17

* Branch 99
Rabr99 node_1 netRa99 484.63340167490566
Lbr99 netRa99 netL99 1.217439918521434e-13
Rbbr99 netL99 node_2 -507.7554862429955
Cbr99 netL99 node_2 5.081285675281899e-19

.ends


* Y'13
.subckt yp13 node_1 node_3
* Branch 0
Rabr0 node_1 netRa0 6100.7944853282925
Lbr0 netRa0 netL0 4.37158519798435e-13
Rbbr0 netL0 node_3 -6121.959115388587
Cbr0 netL0 node_3 1.1743659300624732e-20

* Branch 1
Rabr1 node_1 netRa1 7.624004902960134
Lbr1 netRa1 netL1 -2.5018282605816518e-14
Rbbr1 netL1 node_3 -88.70863696299658
Cbr1 netL1 node_3 -3.245333953686599e-17

* Branch 2
Rabr2 node_1 netRa2 16.20259008922494
Lbr2 netRa2 netL2 -2.4058480468292758e-14
Rbbr2 netL2 node_3 -54.03941238039607
Cbr2 netL2 node_3 -2.589410050595187e-17

* Branch 3
Rabr3 node_1 netRa3 15682.956061987903
Lbr3 netRa3 netL3 1.0268333011441082e-12
Rbbr3 netL3 node_3 -15759.046886735407
Cbr3 netL3 node_3 4.165179492044874e-21

* Branch 4
Rabr4 node_1 netRa4 -4.342330527933723
Lbr4 netRa4 netL4 1.9618851152461113e-14
Rbbr4 netL4 node_3 90.98686737717544
Cbr4 netL4 node_3 4.2825002546102403e-17

* Branch 5
Rabr5 node_1 netRa5 126.63852840824207
Lbr5 netRa5 netL5 6.933072755650766e-14
Rbbr5 netL5 node_3 -241.8935309398391
Cbr5 netL5 node_3 2.3010912412842896e-18

* Branch 6
Rabr6 node_1 netRa6 -42.25913097751124
Lbr6 netRa6 netL6 1.028686662153839e-13
Rbbr6 netL6 node_3 742.2033009708125
Cbr6 netL6 node_3 3.065785280417124e-18

* Branch 7
Rabr7 node_1 netRa7 -5696.465442114616
Lbr7 netRa7 netL7 -1.6378927537888668e-12
Rbbr7 netL7 node_3 6915.968134947506
Cbr7 netL7 node_3 -4.191953521255125e-20

* Branch 8
Rabr8 node_1 netRa8 -29420.25702724363
Lbr8 netRa8 netL8 -5.526007000949021e-12
Rbbr8 netL8 node_3 31814.111349401905
Cbr8 netL8 node_3 -5.935589206482612e-21

* Branch 9
Rabr9 node_1 netRa9 -17069803.11366416
Lbr9 netRa9 netL9 -1.3093064277468318e-10
Rbbr9 netL9 node_3 17072290.74972701
Cbr9 netL9 node_3 -4.493795184666043e-25

* Branch 10
Rabr10 node_1 netRa10 -32670.583656709914
Lbr10 netRa10 netL10 -5.9212454781920995e-12
Rbbr10 netL10 node_3 35221.92861316124
Cbr10 netL10 node_3 -5.171451836124537e-21

* Branch 11
Rabr11 node_1 netRa11 -36.80646706948584
Lbr11 netRa11 netL11 3.574181982018236e-14
Rbbr11 netL11 node_3 52.295066710911144
Cbr11 netL11 node_3 1.8129281666709078e-17

* Branch 12
Rabr12 node_1 netRa12 -1320.850007576878
Lbr12 netRa12 netL12 -3.7776928750672787e-13
Rbbr12 netL12 node_3 1642.5176892370912
Cbr12 netL12 node_3 -1.7537250177476788e-19

* Branch 13
Rabr13 node_1 netRa13 8812.02294224242
Lbr13 netRa13 netL13 -3.1203455029308216e-12
Rbbr13 netL13 node_3 -12476.409155134403
Cbr13 netL13 node_3 -2.8139745283067364e-20

* Branch 14
Rabr14 node_1 netRa14 2416.4979309621995
Lbr14 netRa14 netL14 -1.783170427417568e-12
Rbbr14 netL14 node_3 -6635.295497038413
Cbr14 netL14 node_3 -1.0935626116741855e-19

* Branch 15
Rabr15 node_1 netRa15 -159577.5963282365
Lbr15 netRa15 netL15 1.8598621386622937e-11
Rbbr15 netL15 node_3 164369.15141194814
Cbr15 netL15 node_3 7.071980219365806e-22

* Branch 16
Rabr16 node_1 netRa16 1210.1043579638401
Lbr16 netRa16 netL16 2.43915099148007e-13
Rbbr16 netL16 node_3 -1358.8077442982412
Cbr16 netL16 node_3 1.4901517776549354e-19

* Branch 17
Rabr17 node_1 netRa17 -27556.905202798123
Lbr17 netRa17 netL17 4.816300545380427e-12
Rbbr17 netL17 node_3 29899.184649535193
Cbr17 netL17 node_3 5.824143927594632e-21

* Branch 18
Rabr18 node_1 netRa18 335.45644291601553
Lbr18 netRa18 netL18 -7.099560044757764e-13
Rbbr18 netL18 node_3 -3184.350417536448
Cbr18 netL18 node_3 -6.376547124780636e-19

* Branch 19
Rabr19 node_1 netRa19 956.3911666098548
Lbr19 netRa19 netL19 4.3588744020355214e-13
Rbbr19 netL19 node_3 -1168.3543308627309
Cbr19 netL19 node_3 3.935592502634254e-19

* Branch 20
Rabr20 node_1 netRa20 1267.0503305159277
Lbr20 netRa20 netL20 -8.816682500108051e-13
Rbbr20 netL20 node_3 -3120.846116233018
Cbr20 netL20 node_3 -2.200094323310951e-19

* Branch 21
Rabr21 node_1 netRa21 -263.96837229790754
Lbr21 netRa21 netL21 -8.780092364292501e-13
Rbbr21 netL21 node_3 5673.763769875191
Cbr21 netL21 node_3 -6.252778200041967e-19

* Branch 22
Rabr22 node_1 netRa22 23874992.91785196
Lbr22 netRa22 netL22 -1.778295764193953e-10
Rbbr22 netL22 node_3 -23876261.69522796
Cbr22 netL22 node_3 -3.119132497197715e-25

* Branch 23
Rabr23 node_1 netRa23 24.053212420889075
Lbr23 netRa23 netL23 -4.561583593766815e-13
Rbbr23 netL23 node_3 -13351.424835414635
Cbr23 netL23 node_3 -1.080606275262211e-18

* Branch 24
Rabr24 node_1 netRa24 -56.80445944668897
Lbr24 netRa24 netL24 1.8813600889517472e-13
Rbbr24 netL24 node_3 708.6405927779417
Cbr24 netL24 node_3 4.433424083208929e-18

* Branch 25
Rabr25 node_1 netRa25 -7718.954562761047
Lbr25 netRa25 netL25 -4.169185379397289e-12
Rbbr25 netL25 node_3 13954.001469133438
Cbr25 netL25 node_3 -3.904671026578468e-20

* Branch 26
Rabr26 node_1 netRa26 -758.2047878257405
Lbr26 netRa26 netL26 -1.3154484580444677e-12
Rbbr26 netL26 node_3 4942.308086408788
Cbr26 netL26 node_3 -3.6111257456582e-19

* Branch 27
Rabr27 node_1 netRa27 4708.479868108313
Lbr27 netRa27 netL27 -2.3355419266107144e-12
Rbbr27 netL27 node_3 -6938.912445609109
Cbr27 netL27 node_3 -7.093368631413092e-20

* Branch 28
Rabr28 node_1 netRa28 -72917.49149605485
Lbr28 netRa28 netL28 2.1604332624812618e-12
Rbbr28 netL28 node_3 73050.95701717291
Cbr28 netL28 node_3 4.053998325159935e-22

* Branch 29
Rabr29 node_1 netRa29 45.46472816898843
Lbr29 netRa29 netL29 -2.1754132818437062e-13
Rbbr29 netL29 node_3 -1155.0763116244548
Cbr29 netL29 node_3 -3.8638959614638285e-18

* Branch 30
Rabr30 node_1 netRa30 -0.8250270811652406
Lbr30 netRa30 netL30 1.7471727290929042e-14
Rbbr30 netL30 node_3 125.01338471697566
Cbr30 netL30 node_3 1.2908907600286303e-16

* Branch 31
Rabr31 node_1 netRa31 2583.3342972931227
Lbr31 netRa31 netL31 -4.0975611299371e-12
Rbbr31 netL31 node_3 -18138.600035982483
Cbr31 netL31 node_3 -8.548836296410462e-20

* Branch 32
Rabr32 node_1 netRa32 107.443943448996
Lbr32 netRa32 netL32 -6.400155135336694e-13
Rbbr32 netL32 node_3 -3214.255384757344
Cbr32 netL32 node_3 -1.7081577857413745e-18

* Branch 33
Rabr33 node_1 netRa33 -54350.08548992272
Lbr33 netRa33 netL33 -2.5239528863334e-11
Rbbr33 netL33 node_3 68621.67054409957
Cbr33 netL33 node_3 -6.81196273650896e-21

* Branch 34
Rabr34 node_1 netRa34 260.52186473498784
Lbr34 netRa34 netL34 -1.7353670350880167e-12
Rbbr34 netL34 node_3 -36634.98328172783
Cbr34 netL34 node_3 -1.6621986890727782e-19

* Branch 35
Rabr35 node_1 netRa35 -753.3719193378311
Lbr35 netRa35 netL35 3.1646090365883553e-12
Rbbr35 netL35 node_3 33513.64022125199
Cbr35 netL35 node_3 1.1835799887900862e-19

* Branch 36
Rabr36 node_1 netRa36 1837.8629550099672
Lbr36 netRa36 netL36 -2.1235196112370378e-12
Rbbr36 netL36 node_3 -9584.272455478236
Cbr36 netL36 node_3 -1.186644249723656e-19

* Branch 37
Rabr37 node_1 netRa37 -7654.0780450676675
Lbr37 netRa37 netL37 5.999295857365841e-12
Rbbr37 netL37 node_3 17716.622077040545
Cbr37 netL37 node_3 4.3773753595601734e-20

* Branch 38
Rabr38 node_1 netRa38 -249978.83881342117
Lbr38 netRa38 netL38 -2.7754591222209527e-11
Rbbr38 netL38 node_3 258863.20016267928
Cbr38 netL38 node_3 -4.29543278834037e-22

* Branch 39
Rabr39 node_1 netRa39 4572.039258078593
Lbr39 netRa39 netL39 1.6327469276294369e-12
Rbbr39 netL39 node_3 -5493.256485542332
Cbr39 netL39 node_3 6.531732301124926e-20

* Branch 40
Rabr40 node_1 netRa40 -5237.833315459778
Lbr40 netRa40 netL40 9.88002861777321e-12
Rbbr40 netL40 node_3 67049.23258083062
Cbr40 netL40 node_3 2.7453277931780285e-20

* Branch 41
Rabr41 node_1 netRa41 -16933.759174811854
Lbr41 netRa41 netL41 -3.4607738715105016e-12
Rbbr41 netL41 node_3 17895.18753718323
Cbr41 netL41 node_3 -1.1450107143662728e-20

* Branch 42
Rabr42 node_1 netRa42 18893.489501155695
Lbr42 netRa42 netL42 1.378568146920047e-12
Rbbr42 netL42 node_3 -19102.032752526608
Cbr42 netL42 node_3 3.823112670938334e-21

* Branch 43
Rabr43 node_1 netRa43 6658.761999136487
Lbr43 netRa43 netL43 5.550061292852256e-12
Rbbr43 netL43 node_3 -13069.799836933882
Cbr43 netL43 node_3 6.435922950391476e-20

* Branch 44
Rabr44 node_1 netRa44 43669.434456878145
Lbr44 netRa44 netL44 -2.0755624276043824e-11
Rbbr44 netL44 node_3 -55881.312417246765
Cbr44 netL44 node_3 -8.4616510046087e-21

* Branch 45
Rabr45 node_1 netRa45 -5689.75232336523
Lbr45 netRa45 netL45 -2.5137081377133754e-12
Rbbr45 netL45 node_3 7541.524056162178
Cbr45 netL45 node_3 -5.884828618888738e-20

* Branch 46
Rabr46 node_1 netRa46 -21810.024950723047
Lbr46 netRa46 netL46 9.017832428018755e-12
Rbbr46 netL46 node_3 32352.013085016868
Cbr46 netL46 node_3 1.2727381326823435e-20

* Branch 47
Rabr47 node_1 netRa47 544833.5256696588
Lbr47 netRa47 netL47 -4.874341868700572e-11
Rbbr47 netL47 node_3 -551132.8520209206
Cbr47 netL47 node_3 -1.6218306804244404e-22

* Branch 48
Rabr48 node_1 netRa48 146001.001363157
Lbr48 netRa48 netL48 -2.6460906208390753e-11
Rbbr48 netL48 node_3 -153338.05003485671
Cbr48 netL48 node_3 -1.1798318921621286e-21

* Branch 49
Rabr49 node_1 netRa49 36133.98720797735
Lbr49 netRa49 netL49 1.5871272374949042e-11
Rbbr49 netL49 node_3 -52831.206831785756
Cbr49 netL49 node_3 8.348479949245352e-21

* Branch 50
Rabr50 node_1 netRa50 -38.95983638572261
Lbr50 netRa50 netL50 4.498690282665177e-13
Rbbr50 netL50 node_3 4936.678385846337
Cbr50 netL50 node_3 2.1245519299512915e-18

* Branch 51
Rabr51 node_1 netRa51 -5183.470066244396
Lbr51 netRa51 netL51 -4.1210666314034535e-12
Rbbr51 netL51 node_3 8161.089151253691
Cbr51 netL51 node_3 -9.807756913768407e-20

* Branch 52
Rabr52 node_1 netRa52 206257.2535012941
Lbr52 netRa52 netL52 -1.642147683410019e-11
Rbbr52 netL52 node_3 -207391.1648191749
Cbr52 netL52 node_3 -3.8365889450545134e-22

* Branch 53
Rabr53 node_1 netRa53 53271.97005781572
Lbr53 netRa53 netL53 -1.2548851937701438e-11
Rbbr53 netL53 node_3 -62462.228968308176
Cbr53 netL53 node_3 -3.765189098593202e-21

* Branch 54
Rabr54 node_1 netRa54 -32514.048906531603
Lbr54 netRa54 netL54 -1.1733418838630004e-11
Rbbr54 netL54 node_3 40191.44112066945
Cbr54 netL54 node_3 -8.99896795008342e-21

* Branch 55
Rabr55 node_1 netRa55 9877.775092720081
Lbr55 netRa55 netL55 2.88619881047395e-12
Rbbr55 netL55 node_3 -11662.370391685454
Cbr55 netL55 node_3 2.5099377082357707e-20

* Branch 56
Rabr56 node_1 netRa56 -123235.24238012721
Lbr56 netRa56 netL56 1.7124495337560506e-11
Rbbr56 netL56 node_3 129573.45582131915
Cbr56 netL56 node_3 1.0715501764303305e-21

* Branch 57
Rabr57 node_1 netRa57 580.6820551796504
Lbr57 netRa57 netL57 -3.170650220331964e-12
Rbbr57 netL57 node_3 -22511.692197810407
Cbr57 netL57 node_3 -2.350558875142089e-19

* Branch 58
Rabr58 node_1 netRa58 -2405.78088018367
Lbr58 netRa58 netL58 -8.646463434095623e-12
Rbbr58 netL58 node_3 61053.35825333217
Cbr58 netL58 node_3 -6.011868585473798e-20

* Branch 59
Rabr59 node_1 netRa59 -2004.6223320894612
Lbr59 netRa59 netL59 -4.1129335306224584e-12
Rbbr59 netL59 node_3 18087.300510919325
Cbr59 netL59 node_3 -1.1476473365104453e-19

* Branch 60
Rabr60 node_1 netRa60 -506.4658284936824
Lbr60 netRa60 netL60 -2.2786254751818877e-13
Rbbr60 netL60 node_3 672.7652438982867
Cbr60 netL60 node_3 -6.703513842597324e-19

* Branch 61
Rabr61 node_1 netRa61 5298.908096905543
Lbr61 netRa61 netL61 -6.183578747549649e-12
Rbbr61 netL61 node_3 -14467.91249445974
Cbr61 netL61 node_3 -8.016255588661445e-20

* Branch 62
Rabr62 node_1 netRa62 -1570.5834583685396
Lbr62 netRa62 netL62 4.1162831848559476e-12
Rbbr62 netL62 node_3 12198.57371276208
Cbr62 netL62 node_3 2.1218660675644542e-19

* Branch 63
Rabr63 node_1 netRa63 25553286.634931915
Lbr63 netRa63 netL63 -3.669202976316557e-10
Rbbr63 netL63 node_3 -25566783.292446885
Cbr63 netL63 node_3 -5.61591609996094e-25

* Branch 64
Rabr64 node_1 netRa64 740.0128363298346
Lbr64 netRa64 netL64 -2.7275468635458744e-12
Rbbr64 netL64 node_3 -14017.554141953511
Cbr64 netL64 node_3 -2.593807731116305e-19

* Branch 65
Rabr65 node_1 netRa65 -488.41356337794565
Lbr65 netRa65 netL65 -1.0516816464507443e-12
Rbbr65 netL65 node_3 2376.951996123593
Cbr65 netL65 node_3 -9.112350156083636e-19

* Branch 66
Rabr66 node_1 netRa66 80634.59884034541
Lbr66 netRa66 netL66 -1.4725457829138683e-11
Rbbr66 netL66 node_3 -85242.8156179815
Cbr66 netL66 node_3 -2.1414074092600132e-21

* Branch 67
Rabr67 node_1 netRa67 11336.622334370133
Lbr67 netRa67 netL67 -2.81550200085339e-12
Rbbr67 netL67 node_3 -12454.075591797819
Cbr67 netL67 node_3 -1.9932416470612034e-20

* Branch 68
Rabr68 node_1 netRa68 28376.92548811835
Lbr68 netRa68 netL68 1.7747439262027106e-11
Rbbr68 netL68 node_3 -58260.157571251846
Cbr68 netL68 node_3 1.0746501156956285e-20

* Branch 69
Rabr69 node_1 netRa69 -2441.728761163592
Lbr69 netRa69 netL69 -1.7354489440103834e-12
Rbbr69 netL69 node_3 5002.861952768365
Cbr69 netL69 node_3 -1.4220735364040694e-19

* Branch 70
Rabr70 node_1 netRa70 7231.372586260887
Lbr70 netRa70 netL70 8.682634571884832e-13
Rbbr70 netL70 node_3 -7399.737265437112
Cbr70 netL70 node_3 1.622801408643723e-20

* Branch 71
Rabr71 node_1 netRa71 4729.657674911888
Lbr71 netRa71 netL71 -5.569729462502179e-12
Rbbr71 netL71 node_3 -14404.61740165386
Cbr71 netL71 node_3 -8.16589749432702e-20

* Branch 72
Rabr72 node_1 netRa72 -12617.518421935067
Lbr72 netRa72 netL72 1.9045621690827802e-11
Rbbr72 netL72 node_3 41893.74501835537
Cbr72 netL72 node_3 3.599406866274695e-20

* Branch 73
Rabr73 node_1 netRa73 -922.9624604147788
Lbr73 netRa73 netL73 -7.320368821629329e-12
Rbbr73 netL73 node_3 184655.9733109624
Cbr73 netL73 node_3 -4.3159621153028244e-20

* Branch 74
Rabr74 node_1 netRa74 -1442.0756659850965
Lbr74 netRa74 netL74 -2.1011634997421187e-12
Rbbr74 netL74 node_3 3856.1702740332053
Cbr74 netL74 node_3 -3.7817635713208004e-19

* Branch 75
Rabr75 node_1 netRa75 1911.3326462673847
Lbr75 netRa75 netL75 -4.600091605915114e-12
Rbbr75 netL75 node_3 -18026.442261058608
Cbr75 netL75 node_3 -1.3336098259011347e-19

* Branch 76
Rabr76 node_1 netRa76 2.9419641269030143
Lbr76 netRa76 netL76 3.94566243290985e-12
Rbbr76 netL76 node_3 -5311613.137102967
Cbr76 netL76 node_3 4.793428654940111e-19

* Branch 77
Rabr77 node_1 netRa77 -376.27639239560096
Lbr77 netRa77 netL77 2.970713480954726e-12
Rbbr77 netL77 node_3 12293.982553193517
Cbr77 netL77 node_3 6.40500301394e-19

* Branch 78
Rabr78 node_1 netRa78 982.3080998191185
Lbr78 netRa78 netL78 6.082249041227348e-12
Rbbr78 netL78 node_3 -21672.066782159854
Cbr78 netL78 node_3 2.862147549812069e-19

* Branch 79
Rabr79 node_1 netRa79 26.962003315404708
Lbr79 netRa79 netL79 -1.0834794936653314e-12
Rbbr79 netL79 node_3 -88222.05467449826
Cbr79 netL79 node_3 -4.507641520560426e-19

* Branch 80
Rabr80 node_1 netRa80 -2981.0942111919476
Lbr80 netRa80 netL80 -3.4001020027989562e-12
Rbbr80 netL80 node_3 5947.639230294066
Cbr80 netL80 node_3 -1.918106763623846e-19

* Branch 81
Rabr81 node_1 netRa81 10614.155610975477
Lbr81 netRa81 netL81 1.2180843654227776e-11
Rbbr81 netL81 node_3 -18561.399943205415
Cbr81 netL81 node_3 6.184133399813358e-20

* Branch 82
Rabr82 node_1 netRa82 -679.0202876165099
Lbr82 netRa82 netL82 2.294253215817951e-12
Rbbr82 netL82 node_3 4480.301104334435
Cbr82 netL82 node_3 7.538299876205718e-19

* Branch 83
Rabr83 node_1 netRa83 428886.6009678917
Lbr83 netRa83 netL83 6.09913035027815e-11
Rbbr83 netL83 node_3 -433993.3148795125
Cbr83 netL83 node_3 3.276772048317403e-22

* Branch 84
Rabr84 node_1 netRa84 -719.8680824947509
Lbr84 netRa84 netL84 4.643028670238776e-13
Rbbr84 netL84 node_3 855.027613478183
Cbr84 netL84 node_3 7.543394202182623e-19

* Branch 85
Rabr85 node_1 netRa85 15337.301915497299
Lbr85 netRa85 netL85 1.1127136022713993e-11
Rbbr85 netL85 node_3 -20258.938220211683
Cbr85 netL85 node_3 3.5814552829515936e-20

* Branch 86
Rabr86 node_1 netRa86 1460.2464009297641
Lbr86 netRa86 netL86 4.1927490631512195e-12
Rbbr86 netL86 node_3 -9060.835735098774
Cbr86 netL86 node_3 3.1715351270993846e-19

* Branch 87
Rabr87 node_1 netRa87 -5489.905499660629
Lbr87 netRa87 netL87 -4.90031524999733e-12
Rbbr87 netL87 node_3 8734.21437878367
Cbr87 netL87 node_3 -1.0222979578584128e-19

* Branch 88
Rabr88 node_1 netRa88 -232.80955728516378
Lbr88 netRa88 netL88 2.9251788866798137e-12
Rbbr88 netL88 node_3 24093.229394149133
Cbr88 netL88 node_3 5.189439590365949e-19

* Branch 89
Rabr89 node_1 netRa89 3689.216221006685
Lbr89 netRa89 netL89 2.8397381357314587e-12
Rbbr89 netL89 node_3 -4720.561987093418
Cbr89 netL89 node_3 1.631149556879105e-19

* Branch 90
Rabr90 node_1 netRa90 -2466.7190498713876
Lbr90 netRa90 netL90 3.833190252423426e-12
Rbbr90 netL90 node_3 6480.497664988805
Cbr90 netL90 node_3 2.396289210562693e-19

* Branch 91
Rabr91 node_1 netRa91 -46869.95456365476
Lbr91 netRa91 netL91 1.5570916849386683e-11
Rbbr91 netL91 node_3 50471.91436002183
Cbr91 netL91 node_3 6.581213619126167e-21

* Branch 92
Rabr92 node_1 netRa92 -25306.71487827097
Lbr92 netRa92 netL92 -1.0475770797896063e-11
Rbbr92 netL92 node_3 28424.139465689965
Cbr92 netL92 node_3 -1.456632867730397e-20

* Branch 93
Rabr93 node_1 netRa93 -849.0592311623888
Lbr93 netRa93 netL93 -1.4093763349612645e-12
Rbbr93 netL93 node_3 2745.50027778808
Cbr93 netL93 node_3 -6.051054172622475e-19

* Branch 94
Rabr94 node_1 netRa94 4073602.2614281685
Lbr94 netRa94 netL94 -2.2749088027279455e-10
Rbbr94 netL94 node_3 -4102540.3725804333
Cbr94 netL94 node_3 -1.3611760171888177e-23

* Branch 95
Rabr95 node_1 netRa95 137316.4761095346
Lbr95 netRa95 netL95 -2.310536755033856e-11
Rbbr95 netL95 node_3 -150546.1063447242
Cbr95 netL95 node_3 -1.1171025680530086e-21

* Branch 96
Rabr96 node_1 netRa96 187200.9649257694
Lbr96 netRa96 netL96 -9.90629598803749e-12
Rbbr96 netL96 node_3 -189091.7567151849
Cbr96 netL96 node_3 -2.797108794102569e-22

* Branch 97
Rabr97 node_1 netRa97 4.168063223321889
Lbr97 netRa97 netL97 -1.2803224781200193e-14
Rbbr97 netL97 node_3 -20.90877964277703
Cbr97 netL97 node_3 -1.410508707216578e-16

* Branch 98
Rabr98 node_1 netRa98 -69.51408973156983
Lbr98 netRa98 netL98 -4.7706867963335104e-14
Rbbr98 netL98 node_3 169.7421876400034
Cbr98 netL98 node_3 -4.1215779595275795e-18

* Branch 99
Rabr99 node_1 netRa99 -440.5594219940009
Lbr99 netRa99 netL99 1.0299212396346333e-13
Rbbr99 netL99 node_3 467.6334958187001
Cbr99 netL99 node_3 4.953136387511427e-19

.ends


* Y'14
.subckt yp14 node_1 node_4
* Branch 0
Rabr0 node_1 netRa0 -4.674440532201781
Lbr0 netRa0 netL0 -1.1925071724995389e-14
Rbbr0 netL0 node_4 29.204140388486657
Cbr0 netL0 node_4 -9.84653612722019e-17

* Branch 1
Rabr1 node_1 netRa1 640.7910118557062
Lbr1 netRa1 netL1 7.273228877076872e-13
Rbbr1 netL1 node_4 -995.691913446946
Cbr1 netL1 node_4 1.1973388116416053e-18

* Branch 2
Rabr2 node_1 netRa2 -16.878889321244348
Lbr2 netRa2 netL2 -5.134426183893977e-15
Rbbr2 netL2 node_4 18.66262538441893
Cbr2 netL2 node_4 -1.650324985496039e-17

* Branch 3
Rabr3 node_1 netRa3 -588.8007734251134
Lbr3 netRa3 netL3 -2.7458157685250672e-14
Rbbr3 netL3 node_4 591.4719355195637
Cbr3 netL3 node_4 -7.898032773701458e-20

* Branch 4
Rabr4 node_1 netRa4 -4.638305662656476
Lbr4 netRa4 netL4 -4.225330725131516e-15
Rbbr4 netL4 node_4 12.916914765826332
Cbr4 netL4 node_4 -7.289929589328464e-17

* Branch 5
Rabr5 node_1 netRa5 14.308232189658735
Lbr5 netRa5 netL5 5.17969848295244e-15
Rbbr5 netL5 node_4 -16.447936926075144
Cbr5 netL5 node_4 2.2284531811086674e-17

* Branch 6
Rabr6 node_1 netRa6 0.20083095498559997
Lbr6 netRa6 netL6 -2.2433907660119746e-15
Rbbr6 netL6 node_4 -21.088218462889927
Cbr6 netL6 node_4 -3.875714766406825e-16

* Branch 7
Rabr7 node_1 netRa7 -5.081778839498085
Lbr7 netRa7 netL7 3.666929736605191e-15
Rbbr7 netL7 node_4 8.01578612299309
Cbr7 netL7 node_4 8.795927348261981e-17

* Branch 8
Rabr8 node_1 netRa8 6.877329195778424
Lbr8 netRa8 netL8 5.1130983060141845e-15
Rbbr8 netL8 node_4 -14.97263752266624
Cbr8 netL8 node_4 5.0878764342791796e-17

* Branch 9
Rabr9 node_1 netRa9 4.1928791916569255
Lbr9 netRa9 netL9 -2.255241031873631e-15
Rbbr9 netL9 node_4 -6.680806165706828
Cbr9 netL9 node_4 -7.916612466287351e-17

* Branch 10
Rabr10 node_1 netRa10 268.7551509282625
Lbr10 netRa10 netL10 -1.7378935812765488e-12
Rbbr10 netL10 node_4 -21489.10931021861
Cbr10 netL10 node_4 -2.557449978072539e-19

* Branch 11
Rabr11 node_1 netRa11 9892.775757587664
Lbr11 netRa11 netL11 -9.831445030096853e-13
Rbbr11 netL11 node_4 -10174.564289998281
Cbr11 netL11 node_4 -9.741140292172903e-21

* Branch 12
Rabr12 node_1 netRa12 2379.677145906972
Lbr12 netRa12 netL12 -1.6752359034069712e-12
Rbbr12 netL12 node_4 -4901.678609926649
Cbr12 netL12 node_4 -1.4095335463939996e-19

* Branch 13
Rabr13 node_1 netRa13 -712.955864888125
Lbr13 netRa13 netL13 2.1493275898582846e-12
Rbbr13 netL13 node_4 20623.698689419663
Cbr13 netL13 node_4 1.3549428579639348e-19

* Branch 14
Rabr14 node_1 netRa14 873.7949225238741
Lbr14 netRa14 netL14 1.0422457973533053e-12
Rbbr14 netL14 node_4 -3357.467201654176
Cbr14 netL14 node_4 3.661597856219289e-19

* Branch 15
Rabr15 node_1 netRa15 -278.3105089786751
Lbr15 netRa15 netL15 -1.1626887867627786e-13
Rbbr15 netL15 node_4 381.9105889731116
Cbr15 netL15 node_4 -1.1049211322880726e-18

* Branch 16
Rabr16 node_1 netRa16 20664.410996881026
Lbr16 netRa16 netL16 -4.57158622438203e-12
Rbbr16 netL16 node_4 -23391.554484163353
Cbr16 netL16 node_4 -9.410145605138725e-21

* Branch 17
Rabr17 node_1 netRa17 103.52015756822475
Lbr17 netRa17 netL17 3.792625371160276e-12
Rbbr17 netL17 node_4 -1849775.197381862
Cbr17 netL17 node_4 1.1401713177892219e-19

* Branch 18
Rabr18 node_1 netRa18 250.13418221418905
Lbr18 netRa18 netL18 -3.654104489076378e-13
Rbbr18 netL18 node_4 -476.375793370802
Cbr18 netL18 node_4 -2.971295253463922e-18

* Branch 19
Rabr19 node_1 netRa19 2217.123853891007
Lbr19 netRa19 netL19 1.4961634542684292e-12
Rbbr19 netL19 node_4 -4247.5360751498865
Cbr19 netL19 node_4 1.6122965574577863e-19

* Branch 20
Rabr20 node_1 netRa20 17278.658983295714
Lbr20 netRa20 netL20 6.003376306519108e-12
Rbbr20 netL20 node_4 -22698.024707327953
Cbr20 netL20 node_4 1.5420323042750657e-20

* Branch 21
Rabr21 node_1 netRa21 96101.06757993247
Lbr21 netRa21 netL21 1.2950270589625679e-11
Rbbr21 netL21 node_4 -100313.39380907724
Cbr21 netL21 node_4 1.347045698902163e-21

* Branch 22
Rabr22 node_1 netRa22 -301.5137473807243
Lbr22 netRa22 netL22 2.501542367932836e-13
Rbbr22 netL22 node_4 624.7328512076982
Cbr22 netL22 node_4 1.3062513565060878e-18

* Branch 23
Rabr23 node_1 netRa23 1399.0212908193037
Lbr23 netRa23 netL23 8.172540773824285e-13
Rbbr23 netL23 node_4 -1982.512949109594
Cbr23 netL23 node_4 2.980768518925742e-19

* Branch 24
Rabr24 node_1 netRa24 -465.50387361452727
Lbr24 netRa24 netL24 -1.7122256263293244e-13
Rbbr24 netL24 node_4 595.8765195610401
Cbr24 netL24 node_4 -6.21740166934123e-19

* Branch 25
Rabr25 node_1 netRa25 0.4533882309058711
Lbr25 netRa25 netL25 -2.1742826329426675e-15
Rbbr25 netL25 node_4 -29.095434807685937
Cbr25 netL25 node_4 -1.5147074821005334e-16

* Branch 26
Rabr26 node_1 netRa26 9280.907483266243
Lbr26 netRa26 netL26 1.2387467095716202e-11
Rbbr26 netL26 node_4 -50669.892323613436
Cbr26 netL26 node_4 2.6975681298964808e-20

* Branch 27
Rabr27 node_1 netRa27 233.9989946949526
Lbr27 netRa27 netL27 3.191653607423731e-13
Rbbr27 netL27 node_4 -1602.8630953501104
Cbr27 netL27 node_4 8.718167011967116e-19

* Branch 28
Rabr28 node_1 netRa28 1160.0378689483846
Lbr28 netRa28 netL28 2.291834183977696e-12
Rbbr28 netL28 node_4 -14377.169784089314
Cbr28 netL28 node_4 1.4219847794516267e-19

* Branch 29
Rabr29 node_1 netRa29 1403.0055501811523
Lbr29 netRa29 netL29 2.2873069069708737e-12
Rbbr29 netL29 node_4 -13817.803329578472
Cbr29 netL29 node_4 1.2135151963199346e-19

* Branch 30
Rabr30 node_1 netRa30 12145.649121928856
Lbr30 netRa30 netL30 9.287639246707203e-12
Rbbr30 netL30 node_4 -31038.282434051478
Cbr30 netL30 node_4 2.4956215830076843e-20

* Branch 31
Rabr31 node_1 netRa31 1584.6238352841299
Lbr31 netRa31 netL31 1.1484136118208987e-12
Rbbr31 netL31 node_4 -2629.7959551576614
Cbr31 netL31 node_4 2.7888543976274697e-19

* Branch 32
Rabr32 node_1 netRa32 -637.8560001528685
Lbr32 netRa32 netL32 1.3741084865047065e-12
Rbbr32 netL32 node_4 3209.7250646003085
Cbr32 netL32 node_4 6.483911989001998e-19

* Branch 33
Rabr33 node_1 netRa33 7415.885259289623
Lbr33 netRa33 netL33 1.2261925437799943e-12
Rbbr33 netL33 node_4 -7783.097205063241
Cbr33 netL33 node_4 2.13015525998304e-20

* Branch 34
Rabr34 node_1 netRa34 2663.7926495718852
Lbr34 netRa34 netL34 2.2503603756630316e-12
Rbbr34 netL34 node_4 -5968.286441741068
Cbr34 netL34 node_4 1.4337369140021448e-19

* Branch 35
Rabr35 node_1 netRa35 32.769244048264845
Lbr35 netRa35 netL35 7.15256237984054e-15
Rbbr35 netL35 node_4 -37.46529942759728
Cbr35 netL35 node_4 5.84510804715735e-18

* Branch 36
Rabr36 node_1 netRa36 -3856.2445063810123
Lbr36 netRa36 netL36 1.941886664931217e-12
Rbbr36 netL36 node_4 5351.05262153988
Cbr36 netL36 node_4 9.340525538683832e-20

* Branch 37
Rabr37 node_1 netRa37 -4016.7938684487804
Lbr37 netRa37 netL37 1.2240913118238233e-12
Rbbr37 netL37 node_4 5086.948780337631
Cbr37 netL37 node_4 5.963892769299079e-20

* Branch 38
Rabr38 node_1 netRa38 4107.316871131479
Lbr38 netRa38 netL38 4.338188660365653e-12
Rbbr38 netL38 node_4 -15754.963514930327
Cbr38 netL38 node_4 6.809965061922432e-20

* Branch 39
Rabr39 node_1 netRa39 -26148.19572123003
Lbr39 netRa39 netL39 -6.789226103620444e-12
Rbbr39 netL39 node_4 27817.3563780905
Cbr39 netL39 node_4 -9.369378184821503e-21

* Branch 40
Rabr40 node_1 netRa40 -59498.32115215213
Lbr40 netRa40 netL40 -3.9018256418681725e-11
Rbbr40 netL40 node_4 130413.62771627319
Cbr40 netL40 node_4 -5.07506064455287e-21

* Branch 41
Rabr41 node_1 netRa41 1352.9024601468977
Lbr41 netRa41 netL41 -2.484110858109286e-13
Rbbr41 netL41 node_4 -1404.6090701350154
Cbr41 netL41 node_4 -1.3039032407287123e-19

* Branch 42
Rabr42 node_1 netRa42 -610.2929981508086
Lbr42 netRa42 netL42 3.671876861200944e-12
Rbbr42 netL42 node_4 49054.153166855685
Cbr42 netL42 node_4 1.133370510516243e-19

* Branch 43
Rabr43 node_1 netRa43 -24.53307485687442
Lbr43 netRa43 netL43 5.170486523551693e-15
Rbbr43 netL43 node_4 27.780453763744866
Cbr43 netL43 node_4 7.565157121195753e-18

* Branch 44
Rabr44 node_1 netRa44 -43.816384007048654
Lbr44 netRa44 netL44 3.044299279265799e-13
Rbbr44 netL44 node_4 2172.4899976614215
Cbr44 netL44 node_4 2.9386800833771498e-18

* Branch 45
Rabr45 node_1 netRa45 40367.21197694037
Lbr45 netRa45 netL45 -1.0326148147659395e-11
Rbbr45 netL45 node_4 -43132.63629039442
Cbr45 netL45 node_4 -5.912234386652337e-21

* Branch 46
Rabr46 node_1 netRa46 -235630.50974529446
Lbr46 netRa46 netL46 2.1065286517448707e-11
Rbbr46 netL46 node_4 241993.56052050143
Cbr46 netL46 node_4 3.690341604247065e-22

* Branch 47
Rabr47 node_1 netRa47 284.04050404015675
Lbr47 netRa47 netL47 -7.073216222526764e-13
Rbbr47 netL47 node_4 -3122.091088559238
Cbr47 netL47 node_4 -7.746441401669724e-19

* Branch 48
Rabr48 node_1 netRa48 1323.5383155001396
Lbr48 netRa48 netL48 4.126859076456808e-13
Rbbr48 netL48 node_4 -1497.808264991711
Cbr48 netL48 node_4 2.0891605717835874e-19

* Branch 49
Rabr49 node_1 netRa49 2335.0973231291127
Lbr49 netRa49 netL49 1.5497545802893965e-12
Rbbr49 netL49 node_4 -5567.06494874902
Cbr49 netL49 node_4 1.2010019775630071e-19

* Branch 50
Rabr50 node_1 netRa50 1922.4126370392678
Lbr50 netRa50 netL50 2.2929329702668197e-12
Rbbr50 netL50 node_4 -11437.35350617441
Cbr50 netL50 node_4 1.05682986992698e-19

* Branch 51
Rabr51 node_1 netRa51 -8871.502800311102
Lbr51 netRa51 netL51 3.9847746709868085e-12
Rbbr51 netL51 node_4 10586.579306253027
Cbr51 netL51 node_4 4.2218397806221616e-20

* Branch 52
Rabr52 node_1 netRa52 -363.72696752535387
Lbr52 netRa52 netL52 1.1498501845218938e-12
Rbbr52 netL52 node_4 6594.352798887327
Cbr52 netL52 node_4 4.638105361279819e-19

* Branch 53
Rabr53 node_1 netRa53 -5.410843168071725
Lbr53 netRa53 netL53 1.2366141946616008e-12
Rbbr53 netL53 node_4 72843.46571229813
Cbr53 netL53 node_4 9.333928711742426e-19

* Branch 54
Rabr54 node_1 netRa54 116999374005.09827
Lbr54 netRa54 netL54 -1.4347465778424626e-08
Rbbr54 netL54 node_4 -116999377307.864
Cbr54 netL54 node_4 -1.0481116934399299e-30

* Branch 55
Rabr55 node_1 netRa55 21791.55184511536
Lbr55 netRa55 netL55 7.458234573737965e-12
Rbbr55 netL55 node_4 -28632.863044799957
Cbr55 netL55 node_4 1.1994436468099553e-20

* Branch 56
Rabr56 node_1 netRa56 3908.8504593063817
Lbr56 netRa56 netL56 2.1325716582074466e-12
Rbbr56 netL56 node_4 -7642.151135875994
Cbr56 netL56 node_4 7.177878690119826e-20

* Branch 57
Rabr57 node_1 netRa57 112.3521658250491
Lbr57 netRa57 netL57 -6.563690166527926e-13
Rbbr57 netL57 node_4 -5086.9191534456695
Cbr57 netL57 node_4 -1.0874338315220164e-18

* Branch 58
Rabr58 node_1 netRa58 7114.523264601568
Lbr58 netRa58 netL58 5.417352461998659e-13
Rbbr58 netL58 node_4 -7181.364649568854
Cbr58 netL58 node_4 1.0610840409866368e-20

* Branch 59
Rabr59 node_1 netRa59 868.5271997834826
Lbr59 netRa59 netL59 1.4899569384384129e-12
Rbbr59 netL59 node_4 -4583.523799904036
Cbr59 netL59 node_4 3.803712687416445e-19

* Branch 60
Rabr60 node_1 netRa60 42696.98757045408
Lbr60 netRa60 netL60 1.3153646579758932e-11
Rbbr60 netL60 node_4 -52986.78911845618
Cbr60 netL60 node_4 5.827988956345642e-21

* Branch 61
Rabr61 node_1 netRa61 -601.0306725372706
Lbr61 netRa61 netL61 1.172980822509305e-12
Rbbr61 netL61 node_4 3489.868186280467
Cbr61 netL61 node_4 5.510532705679997e-19

* Branch 62
Rabr62 node_1 netRa62 -53.722857613892145
Lbr62 netRa62 netL62 5.99410781250577e-13
Rbbr62 netL62 node_4 8122.711471196811
Cbr62 netL62 node_4 1.2664101137676566e-18

* Branch 63
Rabr63 node_1 netRa63 -71753.74358733988
Lbr63 netRa63 netL63 2.381154469759006e-11
Rbbr63 netL63 node_4 79783.11327485576
Cbr63 netL63 node_4 4.150871547048939e-21

* Branch 64
Rabr64 node_1 netRa64 8214.283411516488
Lbr64 netRa64 netL64 -2.4300567186964624e-12
Rbbr64 netL64 node_4 -8810.368614846593
Cbr64 netL64 node_4 -3.351726683258176e-20

* Branch 65
Rabr65 node_1 netRa65 36279.74758759918
Lbr65 netRa65 netL65 1.0368135608105692e-11
Rbbr65 netL65 node_4 -40649.42951856917
Cbr65 netL65 node_4 7.041065956950885e-21

* Branch 66
Rabr66 node_1 netRa66 -101006.69138945667
Lbr66 netRa66 netL66 9.263891874941802e-12
Rbbr66 netL66 node_4 102542.24097680338
Cbr66 netL66 node_4 8.940258946308503e-22

* Branch 67
Rabr67 node_1 netRa67 -554.9885170306945
Lbr67 netRa67 netL67 6.993913557581069e-13
Rbbr67 netL67 node_4 1729.9187794827387
Cbr67 netL67 node_4 7.250881474396228e-19

* Branch 68
Rabr68 node_1 netRa68 381.59166532738465
Lbr68 netRa68 netL68 -8.044191665650959e-14
Rbbr68 netL68 node_4 -394.91863921837825
Cbr68 netL68 node_4 -5.334151500675209e-19

* Branch 69
Rabr69 node_1 netRa69 -6285.6425610956285
Lbr69 netRa69 netL69 -6.450778445841449e-12
Rbbr69 netL69 node_4 12898.338867754128
Cbr69 netL69 node_4 -7.984118961983629e-20

* Branch 70
Rabr70 node_1 netRa70 4368.264720990602
Lbr70 netRa70 netL70 2.7915013921568503e-12
Rbbr70 netL70 node_4 -6959.657429459465
Cbr70 netL70 node_4 9.193580961853964e-20

* Branch 71
Rabr71 node_1 netRa71 8160260.35166237
Lbr71 netRa71 netL71 2.5430326698890673e-10
Rbbr71 netL71 node_4 -8185260.570433365
Cbr71 netL71 node_4 3.80743981136153e-24

* Branch 72
Rabr72 node_1 netRa72 -170.56624323560877
Lbr72 netRa72 netL72 -1.701370207051555e-13
Rbbr72 netL72 node_4 444.2054273738833
Cbr72 netL72 node_4 -2.2479552446709043e-18

* Branch 73
Rabr73 node_1 netRa73 -77869.75331573824
Lbr73 netRa73 netL73 -2.2968124870114335e-11
Rbbr73 netL73 node_4 93446.46918596652
Cbr73 netL73 node_4 -3.1573443944633413e-21

* Branch 74
Rabr74 node_1 netRa74 -319.0944586746403
Lbr74 netRa74 netL74 -3.814058649179928e-12
Rbbr74 netL74 node_4 23781.039395409258
Cbr74 netL74 node_4 -5.078749520478057e-19

* Branch 75
Rabr75 node_1 netRa75 -191.89309533265902
Lbr75 netRa75 netL75 -3.5331113801032303e-12
Rbbr75 netL75 node_4 32584.95704443417
Cbr75 netL75 node_4 -5.735981699993012e-19

* Branch 76
Rabr76 node_1 netRa76 -450.9607728797192
Lbr76 netRa76 netL76 -4.217945510240525e-12
Rbbr76 netL76 node_4 21446.898272039653
Cbr76 netL76 node_4 -4.391326626253058e-19

* Branch 77
Rabr77 node_1 netRa77 -487.0366829618211
Lbr77 netRa77 netL77 -5.573245299689348e-12
Rbbr77 netL77 node_4 35716.147695694635
Cbr77 netL77 node_4 -3.228231749266425e-19

* Branch 78
Rabr78 node_1 netRa78 -573.5518596932269
Lbr78 netRa78 netL78 -6.938802414767543e-12
Rbbr78 netL78 node_4 48599.41118850643
Cbr78 netL78 node_4 -2.506221474486106e-19

* Branch 79
Rabr79 node_1 netRa79 -1439.0656377942598
Lbr79 netRa79 netL79 -8.05967169020991e-12
Rbbr79 netL79 node_4 28060.166356262213
Cbr79 netL79 node_4 -1.999652930991999e-19

* Branch 80
Rabr80 node_1 netRa80 -32.28024837648067
Lbr80 netRa80 netL80 -2.6385267867602883e-12
Rbbr80 netL80 node_4 102247.27279653751
Cbr80 netL80 node_4 -8.028873485281682e-19

* Branch 81
Rabr81 node_1 netRa81 -4366.673625050216
Lbr81 netRa81 netL81 -9.627923359181511e-12
Rbbr81 netL81 node_4 17306.740166098036
Cbr81 netL81 node_4 -1.2741362746438448e-19

* Branch 82
Rabr82 node_1 netRa82 -145.07792290220831
Lbr82 netRa82 netL82 1.3296928342255588e-13
Rbbr82 netL82 node_4 342.76965921640914
Cbr82 netL82 node_4 2.673745724153192e-18

* Branch 83
Rabr83 node_1 netRa83 1254.8694844241356
Lbr83 netRa83 netL83 -7.550689914921813e-12
Rbbr83 netL83 node_4 -29877.560376876547
Cbr83 netL83 node_4 -2.0114183862013943e-19

* Branch 84
Rabr84 node_1 netRa84 26.77013946049782
Lbr84 netRa84 netL84 -1.8783312327631583e-13
Rbbr84 netL84 node_4 -1088.9305780166262
Cbr84 netL84 node_4 -6.430801872609776e-18

* Branch 85
Rabr85 node_1 netRa85 8.406208028861114
Lbr85 netRa85 netL85 2.113459314161545e-13
Rbbr85 netL85 node_4 -4103.810224861508
Cbr85 netL85 node_4 6.174366062128413e-18

* Branch 86
Rabr86 node_1 netRa86 19115.875745871657
Lbr86 netRa86 netL86 -1.1244353772790208e-11
Rbbr86 netL86 node_4 -23430.303645869593
Cbr86 netL86 node_4 -2.5099090466732372e-20

* Branch 87
Rabr87 node_1 netRa87 44044.35066437332
Lbr87 netRa87 netL87 1.179212532059487e-11
Rbbr87 netL87 node_4 -46173.92957581387
Cbr87 netL87 node_4 5.799218199833482e-21

* Branch 88
Rabr88 node_1 netRa88 1708.818326939438
Lbr88 netRa88 netL88 1.664114392678188e-12
Rbbr88 netL88 node_4 -2838.4208377971418
Cbr88 netL88 node_4 3.4332584407722396e-19

* Branch 89
Rabr89 node_1 netRa89 28.666167321316603
Lbr89 netRa89 netL89 3.0640596442846456e-13
Rbbr89 netL89 node_4 -2478.7757419526965
Cbr89 netL89 node_4 4.350190914443398e-18

* Branch 90
Rabr90 node_1 netRa90 12015.773052133078
Lbr90 netRa90 netL90 1.71938868824867e-11
Rbbr90 netL90 node_4 -95772.29374474431
Cbr90 netL90 node_4 1.4959777361676955e-20

* Branch 91
Rabr91 node_1 netRa91 209.11410228828763
Lbr91 netRa91 netL91 4.926241933607197e-13
Rbbr91 netL91 node_4 -1045.087808159015
Cbr91 netL91 node_4 2.258802358898165e-18

* Branch 92
Rabr92 node_1 netRa92 -12.839626005135376
Lbr92 netRa92 netL92 1.5852378193479188e-14
Rbbr92 netL92 node_4 28.166047411759486
Cbr92 netL92 node_4 4.377755527060449e-17

* Branch 93
Rabr93 node_1 netRa93 456.70682788889815
Lbr93 netRa93 netL93 1.2362294749164446e-12
Rbbr93 netL93 node_4 -1977.940523457909
Cbr93 netL93 node_4 1.374222509471901e-18

* Branch 94
Rabr94 node_1 netRa94 11508508.368687894
Lbr94 netRa94 netL94 2.8576275630313085e-10
Rbbr94 netL94 node_4 -11521657.211972997
Cbr94 netL94 node_4 2.155220147684167e-24

* Branch 95
Rabr95 node_1 netRa95 -362766.1660706773
Lbr95 netRa95 netL95 -1.3612653423533984e-11
Rbbr95 netL95 node_4 364608.5906550885
Cbr95 netL95 node_4 -1.0293838584027202e-22

* Branch 96
Rabr96 node_1 netRa96 -87248.35021764929
Lbr96 netRa96 netL96 -6.0466582924106335e-12
Rbbr96 netL96 node_4 87434.12369220592
Cbr96 netL96 node_4 -7.930143064250636e-22

* Branch 97
Rabr97 node_1 netRa97 11.160538018788126
Lbr97 netRa97 netL97 8.281232753751117e-15
Rbbr97 netL97 node_4 -29.666942909371485
Cbr97 netL97 node_4 2.5176873606173597e-17

* Branch 98
Rabr98 node_1 netRa98 -0.03263304877054025
Lbr98 netRa98 netL98 1.8700577073470607e-15
Rbbr98 netL98 node_4 80.00789585656901
Cbr98 netL98 node_4 2.572332032408117e-16

* Branch 99
Rabr99 node_1 netRa99 10.526587182113865
Lbr99 netRa99 netL99 5.144518172750042e-15
Rbbr99 netL99 node_4 -13.440870984963722
Cbr99 netL99 node_4 3.7009053774647466e-17

.ends


* Y'22
.subckt yp22 node_2 0
* Branch 0
Rabr0 node_2 netRa0 367.68060993442145
Lbr0 netRa0 netL0 1.7357440776114356e-12
Rbbr0 netL0 0 -14028.521654352255
Cbr0 netL0 0 3.831257409024969e-19

* Branch 1
Rabr1 node_2 netRa1 1788005.58064676
Lbr1 netRa1 netL1 -6.884331077416979e-10
Rbbr1 netL1 0 -2036935.2597638287
Cbr1 netL1 0 -1.873796496607082e-22

* Branch 2
Rabr2 node_2 netRa2 200938.42437194902
Lbr2 netRa2 netL2 3.198871933423173e-11
Rbbr2 netL2 0 -217309.5018572862
Cbr2 netL2 0 7.352202998446094e-22

* Branch 3
Rabr3 node_2 netRa3 6344.227368076897
Lbr3 netRa3 netL3 4.7014472155194576e-12
Rbbr3 netL3 0 -17410.681010852037
Cbr3 netL3 0 4.3067701017032695e-20

* Branch 4
Rabr4 node_2 netRa4 -247067.00949310782
Lbr4 netRa4 netL4 -2.572341520187361e-11
Rbbr4 netL4 0 251938.93364915022
Cbr4 netL4 0 -4.1385149956972986e-22

* Branch 5
Rabr5 node_2 netRa5 91446.69794286348
Lbr5 netRa5 netL5 2.8579635885086137e-11
Rbbr5 netL5 0 -107766.91459231188
Cbr5 netL5 0 2.9124553577338428e-21

* Branch 6
Rabr6 node_2 netRa6 -1163.5177810732273
Lbr6 netRa6 netL6 2.251175939968205e-12
Rbbr6 netL6 0 14037.260105814552
Cbr6 netL6 0 1.3443053367669398e-19

* Branch 7
Rabr7 node_2 netRa7 -484.4478624986917
Lbr7 netRa7 netL7 -3.2977901026675317e-12
Rbbr7 netL7 0 79999.93794175374
Cbr7 netL7 0 -9.336887215275775e-20

* Branch 8
Rabr8 node_2 netRa8 -92413.9016814756
Lbr8 netRa8 netL8 5.7309521562728575e-11
Rbbr8 netL8 0 184151.83583997842
Cbr8 netL8 0 3.3424872900938813e-21

* Branch 9
Rabr9 node_2 netRa9 18047.983686508636
Lbr9 netRa9 netL9 -2.7331889271986643e-11
Rbbr9 netL9 0 -56361.86704839108
Cbr9 netL9 0 -2.638874435929117e-20

* Branch 10
Rabr10 node_2 netRa10 -20486.471050800876
Lbr10 netRa10 netL10 -8.737695892599126e-12
Rbbr10 netL10 0 28696.954240009236
Cbr10 netL10 0 -1.4924700020492763e-20

* Branch 11
Rabr11 node_2 netRa11 -21924.146809607435
Lbr11 netRa11 netL11 4.902434001849001e-11
Rbbr11 netL11 0 397928.8609511749
Cbr11 netL11 0 5.499557002273496e-21

* Branch 12
Rabr12 node_2 netRa12 -78260.98440256975
Lbr12 netRa12 netL12 -1.3581904525669652e-10
Rbbr12 netL12 0 544103.2049381727
Cbr12 netL12 0 -3.2233350824763863e-21

* Branch 13
Rabr13 node_2 netRa13 1055.333316337117
Lbr13 netRa13 netL13 -9.760809407070928e-12
Rbbr13 netL13 0 -81320.04652405431
Cbr13 netL13 0 -1.0919420128870007e-19

* Branch 14
Rabr14 node_2 netRa14 -4569.025451226142
Lbr14 netRa14 netL14 4.1912778142262325e-12
Rbbr14 netL14 0 6433.810595115176
Cbr14 netL14 0 1.4201697974064706e-19

* Branch 15
Rabr15 node_2 netRa15 207130296.48375475
Lbr15 netRa15 netL15 -2.664547534249028e-09
Rbbr15 netL15 0 -207245064.8314647
Cbr15 netL15 0 -6.206861956945372e-26

* Branch 16
Rabr16 node_2 netRa16 -757512.0037004756
Lbr16 netRa16 netL16 -3.866049273237171e-10
Rbbr16 netL16 0 927172.9589253129
Cbr16 netL16 0 -5.515851095664274e-22

* Branch 17
Rabr17 node_2 netRa17 812808.9544155123
Lbr17 netRa17 netL17 1.6141407531563193e-10
Rbbr17 netL17 0 -862089.3376779357
Cbr17 netL17 0 2.304532512250019e-22

* Branch 18
Rabr18 node_2 netRa18 -2138032.9347568364
Lbr18 netRa18 netL18 1.1807312221229359e-09
Rbbr18 netL18 0 2821063.1352496184
Cbr18 netL18 0 1.9553823047619965e-22

* Branch 19
Rabr19 node_2 netRa19 -316562.0278333906
Lbr19 netRa19 netL19 -3.875412951602801e-10
Rbbr19 netL19 0 691680.4504432521
Cbr19 netL19 0 -1.7740971504989612e-21

* Branch 20
Rabr20 node_2 netRa20 -1395124235.4860406
Lbr20 netRa20 netL20 1.2895566339229324e-08
Rbbr20 netL20 0 1395445712.8675282
Cbr20 netL20 0 6.623806945283092e-27

* Branch 21
Rabr21 node_2 netRa21 1531037.4460641171
Lbr21 netRa21 netL21 -1.068235024831935e-09
Rbbr21 netL21 0 -2288182.7220716313
Cbr21 netL21 0 -3.0459975832175155e-22

* Branch 22
Rabr22 node_2 netRa22 691.9645581954185
Lbr22 netRa22 netL22 -1.4785886733426766e-10
Rbbr22 netL22 0 -52648610.529336736
Cbr22 netL22 0 -3.141665020729987e-21

* Branch 23
Rabr23 node_2 netRa23 -1670177.4104579736
Lbr23 netRa23 netL23 5.612383810185408e-10
Rbbr23 netL23 0 2130000.604267909
Cbr23 netL23 0 1.5769948275529332e-22

* Branch 24
Rabr24 node_2 netRa24 56550.39474477246
Lbr24 netRa24 netL24 -1.0300852126043139e-10
Rbbr24 netL24 0 -141417.53772823914
Cbr24 netL24 0 -1.2852999877309599e-20

* Branch 25
Rabr25 node_2 netRa25 319197.58958503656
Lbr25 netRa25 netL25 1.9762556894662195e-10
Rbbr25 netL25 0 -523816.1340620721
Cbr25 netL25 0 1.1827131274791944e-21

* Branch 26
Rabr26 node_2 netRa26 -1059828.5391015196
Lbr26 netRa26 netL26 -4.612039107494131e-10
Rbbr26 netL26 0 1619510.4511220905
Cbr26 netL26 0 -2.6882114005575833e-22

* Branch 27
Rabr27 node_2 netRa27 -521239.0686743962
Lbr27 netRa27 netL27 -4.579487833597737e-10
Rbbr27 netL27 0 1372808.9848356675
Cbr27 netL27 0 -6.4054649935264605e-22

* Branch 28
Rabr28 node_2 netRa28 -674595.8048117363
Lbr28 netRa28 netL28 -3.1815654336324023e-10
Rbbr28 netL28 0 1106684.093952832
Cbr28 netL28 0 -4.263547356310426e-22

* Branch 29
Rabr29 node_2 netRa29 -1060063.2889313865
Lbr29 netRa29 netL29 1.301041524332724e-09
Rbbr29 netL29 0 2463462.703873088
Cbr29 netL29 0 4.9768162722565245e-22

* Branch 30
Rabr30 node_2 netRa30 327.8477051797903
Lbr30 netRa30 netL30 -4.896481026786274e-11
Rbbr30 netL30 0 -12168552.687275678
Cbr30 netL30 0 -1.0870960509714679e-20

* Branch 31
Rabr31 node_2 netRa31 131229.10426870116
Lbr31 netRa31 netL31 -1.8697645396241218e-10
Rbbr31 netL31 0 -247161.05829526868
Cbr31 netL31 0 -5.757729173318727e-21

* Branch 32
Rabr32 node_2 netRa32 -36277.67413573622
Lbr32 netRa32 netL32 2.0725305304638245e-10
Rbbr32 netL32 0 2811165.704964944
Cbr32 netL32 0 2.02310643119009e-21

* Branch 33
Rabr33 node_2 netRa33 -484090.85391502734
Lbr33 netRa33 netL33 4.481163054681948e-10
Rbbr33 netL33 0 1477736.1037079876
Cbr33 netL33 0 6.260201518382599e-22

* Branch 34
Rabr34 node_2 netRa34 -322732.3038884795
Lbr34 netRa34 netL34 -3.2070401931522826e-10
Rbbr34 netL34 0 1197400.0161628
Cbr34 netL34 0 -8.303911188854566e-22

* Branch 35
Rabr35 node_2 netRa35 48439.07067063246
Lbr35 netRa35 netL35 -1.3167567437833577e-10
Rbbr35 netL35 0 -584806.8053093649
Cbr35 netL35 0 -4.6412112596085434e-21

* Branch 36
Rabr36 node_2 netRa36 2535494.1817035037
Lbr36 netRa36 netL36 8.346249321082696e-10
Rbbr36 netL36 0 -2985019.0451686685
Cbr36 netL36 0 1.1029567453571054e-22

* Branch 37
Rabr37 node_2 netRa37 -79013.33539312656
Lbr37 netRa37 netL37 7.024037212859157e-11
Rbbr37 netL37 0 201969.70326602814
Cbr37 netL37 0 4.399416018287878e-21

* Branch 38
Rabr38 node_2 netRa38 147197.0039278541
Lbr38 netRa38 netL38 -2.424798802998265e-10
Rbbr38 netL38 0 -314039.4717568334
Cbr38 netL38 0 -5.24130865828541e-21

* Branch 39
Rabr39 node_2 netRa39 2099.454122579015
Lbr39 netRa39 netL39 2.947840893792151e-11
Rbbr39 netL39 0 -412533.7659344224
Cbr39 netL39 0 3.425588854245399e-20

* Branch 40
Rabr40 node_2 netRa40 692464.9040186919
Lbr40 netRa40 netL40 1.5463190698421208e-10
Rbbr40 netL40 0 -770659.6801373174
Cbr40 netL40 0 2.897879479016471e-22

* Branch 41
Rabr41 node_2 netRa41 -506865.95380190504
Lbr41 netRa41 netL41 -1.195168279999787e-10
Rbbr41 netL41 0 591861.3074469808
Cbr41 netL41 0 -3.984339743942501e-22

* Branch 42
Rabr42 node_2 netRa42 97190.80085592205
Lbr42 netRa42 netL42 2.7653171848012716e-10
Rbbr42 netL42 0 -1919307.4050007681
Cbr42 netL42 0 1.4839299291919977e-21

* Branch 43
Rabr43 node_2 netRa43 187998.71762393744
Lbr43 netRa43 netL43 -3.184835933151425e-10
Rbbr43 netL43 0 -404071.671739942
Cbr43 netL43 0 -4.190035876269807e-21

* Branch 44
Rabr44 node_2 netRa44 -89251869.50763284
Lbr44 netRa44 netL44 -3.80073563998459e-09
Rbbr44 netL44 0 89732526.04014191
Cbr44 netL44 0 -4.745761462151261e-25

* Branch 45
Rabr45 node_2 netRa45 -82747.47140715363
Lbr45 netRa45 netL45 1.7147443298096554e-10
Rbbr45 netL45 0 270205.3566955017
Cbr45 netL45 0 7.665743287081094e-21

* Branch 46
Rabr46 node_2 netRa46 -3735041.561433093
Lbr46 netRa46 netL46 2.0922925299465645e-09
Rbbr46 netL46 0 6693207.692700097
Cbr46 netL46 0 8.368830946391077e-23

* Branch 47
Rabr47 node_2 netRa47 -26687237.706011716
Lbr47 netRa47 netL47 -3.808555783459534e-09
Rbbr47 netL47 0 27103300.334039167
Cbr47 netL47 0 -5.265520109333957e-24

* Branch 48
Rabr48 node_2 netRa48 -808399.6139975113
Lbr48 netRa48 netL48 8.027934437387968e-10
Rbbr48 netL48 0 1328328.8414194465
Cbr48 netL48 0 7.475453090654412e-22

* Branch 49
Rabr49 node_2 netRa49 -11130041.679149719
Lbr49 netRa49 netL49 2.7947612312510646e-09
Rbbr49 netL49 0 11634309.201901648
Cbr49 netL49 0 2.158239645694792e-23

* Branch 50
Rabr50 node_2 netRa50 769639.8266031435
Lbr50 netRa50 netL50 -1.2972206476846272e-08
Rbbr50 netL50 0 -162994797.8871453
Cbr50 netL50 0 -1.033285633351352e-22

* Branch 51
Rabr51 node_2 netRa51 48013.39292767459
Lbr51 netRa51 netL51 1.70341582350218e-10
Rbbr51 netL51 0 -696673.6149842606
Cbr51 netL51 0 5.092527895740126e-21

* Branch 52
Rabr52 node_2 netRa52 -5561520.278547425
Lbr52 netRa52 netL52 2.5090963776436544e-09
Rbbr52 netL52 0 8370624.2165754335
Cbr52 netL52 0 5.389564058116591e-23

* Branch 53
Rabr53 node_2 netRa53 -7918766.573494217
Lbr53 netRa53 netL53 2.579346049523114e-09
Rbbr53 netL53 0 8485124.264734885
Cbr53 netL53 0 3.8387013858524536e-23

* Branch 54
Rabr54 node_2 netRa54 -275452.9316185723
Lbr54 netRa54 netL54 3.02662078109402e-10
Rbbr54 netL54 0 457523.2219182393
Cbr54 netL54 0 2.4013579221175496e-21

* Branch 55
Rabr55 node_2 netRa55 -448217.1372028119
Lbr55 netRa55 netL55 3.9723099110517823e-10
Rbbr55 netL55 0 1351242.8751992139
Cbr55 netL55 0 6.558074421675609e-22

* Branch 56
Rabr56 node_2 netRa56 63172.26180131325
Lbr56 netRa56 netL56 1.1524634246831777e-09
Rbbr56 netL56 0 -59722778.15643582
Cbr56 netL56 0 3.0612917322703665e-22

* Branch 57
Rabr57 node_2 netRa57 -3562417.1294349055
Lbr57 netRa57 netL57 -2.025200230736733e-09
Rbbr57 netL57 0 4364448.3979248125
Cbr57 netL57 0 -1.3026414739392583e-22

* Branch 58
Rabr58 node_2 netRa58 28203.617433902815
Lbr58 netRa58 netL58 2.613168684361802e-10
Rbbr58 netL58 0 -2838159.033420589
Cbr58 netL58 0 3.2684555157070724e-21

* Branch 59
Rabr59 node_2 netRa59 -46637.83259392415
Lbr59 netRa59 netL59 -5.813844891157754e-10
Rbbr59 netL59 0 4474600.929004054
Cbr59 netL59 0 -2.7914473452970344e-21

* Branch 60
Rabr60 node_2 netRa60 -48060.13105743202
Lbr60 netRa60 netL60 -5.095161308730905e-10
Rbbr60 netL60 0 3234775.2812048183
Cbr60 netL60 0 -3.2831789874788863e-21

* Branch 61
Rabr61 node_2 netRa61 -2178251.4690730427
Lbr61 netRa61 netL61 -1.2848678177328042e-09
Rbbr61 netL61 0 2656370.941464634
Cbr61 netL61 0 -2.2207740348924775e-22

* Branch 62
Rabr62 node_2 netRa62 -6996.228971755374
Lbr62 netRa62 netL62 2.5823746952467315e-10
Rbbr62 netL62 0 10709683.17196652
Cbr62 netL62 0 3.4231535761422866e-21

* Branch 63
Rabr63 node_2 netRa63 -266378.83620361186
Lbr63 netRa63 netL63 1.6700558736030743e-10
Rbbr63 netL63 0 319469.20058956335
Cbr63 netL63 0 1.962197205116974e-21

* Branch 64
Rabr64 node_2 netRa64 -3061500.9717418645
Lbr64 netRa64 netL64 9.08562291030673e-10
Rbbr64 netL64 0 3286535.333946118
Cbr64 netL64 0 9.029230488678728e-23

* Branch 65
Rabr65 node_2 netRa65 55865.13242390456
Lbr65 netRa65 netL65 -1.8957065141061917e-10
Rbbr65 netL65 0 -918098.3052174057
Cbr65 netL65 0 -3.693021095401832e-21

* Branch 66
Rabr66 node_2 netRa66 -321321.22667211393
Lbr66 netRa66 netL66 -4.911407018625376e-10
Rbbr66 netL66 0 748085.617839443
Cbr66 netL66 0 -2.043995829511268e-21

* Branch 67
Rabr67 node_2 netRa67 4638.315774888381
Lbr67 netRa67 netL67 -1.7439744983492236e-10
Rbbr67 netL67 0 -8918443.942879733
Cbr67 netL67 0 -4.175294769317346e-21

* Branch 68
Rabr68 node_2 netRa68 23948.356946656593
Lbr68 netRa68 netL68 -2.367362404048718e-10
Rbbr68 netL68 0 -3082178.6403303896
Cbr68 netL68 0 -3.198774604836458e-21

* Branch 69
Rabr69 node_2 netRa69 -2071.6258131506297
Lbr69 netRa69 netL69 -1.2933120050939855e-10
Rbbr69 netL69 0 11539969.44809891
Cbr69 netL69 0 -5.504794157168167e-21

* Branch 70
Rabr70 node_2 netRa70 -1060546.4929233852
Lbr70 netRa70 netL70 -7.055236109515687e-10
Rbbr70 netL70 0 1618946.1125476565
Cbr70 netL70 0 -4.109968350764647e-22

* Branch 71
Rabr71 node_2 netRa71 -740287.3011897895
Lbr71 netRa71 netL71 6.284257245839098e-10
Rbbr71 netL71 0 1328319.7125970551
Cbr71 netL71 0 6.389053775191374e-22

* Branch 72
Rabr72 node_2 netRa72 1840.5338133417308
Lbr72 netRa72 netL72 -8.306221825295569e-11
Rbbr72 netL72 0 -5305911.745060287
Cbr72 netL72 0 -8.37821627758024e-21

* Branch 73
Rabr73 node_2 netRa73 -10566865.260084813
Lbr73 netRa73 netL73 -2.2964090115351747e-09
Rbbr73 netL73 0 11190218.665406011
Cbr73 netL73 0 -1.94221214810864e-23

* Branch 74
Rabr74 node_2 netRa74 -128943.11857883078
Lbr74 netRa74 netL74 -2.9153630096203806e-10
Rbbr74 netL74 0 972998.527438622
Cbr74 netL74 0 -2.3255216143177865e-21

* Branch 75
Rabr75 node_2 netRa75 -11450.136844314853
Lbr75 netRa75 netL75 4.255437962212735e-11
Rbbr75 netL75 0 472045.2786093135
Cbr75 netL75 0 7.86265172008623e-21

* Branch 76
Rabr76 node_2 netRa76 644894.7892001172
Lbr76 netRa76 netL76 -3.767867892691894e-10
Rbbr76 netL76 0 -990100.2610991643
Cbr76 netL76 0 -5.899760890557463e-22

* Branch 77
Rabr77 node_2 netRa77 -855239.5102914304
Lbr77 netRa77 netL77 -6.489684827677582e-10
Rbbr77 netL77 0 1455795.6607828487
Cbr77 netL77 0 -5.213875930672182e-22

* Branch 78
Rabr78 node_2 netRa78 -176892.39871758834
Lbr78 netRa78 netL78 -1.2958768606967126e-10
Rbbr78 netL78 0 429433.3041100054
Cbr78 netL78 0 -1.7063986776356787e-21

* Branch 79
Rabr79 node_2 netRa79 20191.266443588913
Lbr79 netRa79 netL79 8.758056963994358e-11
Rbbr79 netL79 0 -855033.7619679188
Cbr79 netL79 0 5.081647707084295e-21

* Branch 80
Rabr80 node_2 netRa80 25641.350539327508
Lbr80 netRa80 netL80 1.7091163401454135e-10
Rbbr80 netL80 0 -2577934.773448138
Cbr80 netL80 0 2.593700104914631e-21

* Branch 81
Rabr81 node_2 netRa81 108085.99165767491
Lbr81 netRa81 netL81 -1.1989656529067408e-10
Rbbr81 netL81 0 -344506.75594781036
Cbr81 netL81 0 -3.218010839195713e-21

* Branch 82
Rabr82 node_2 netRa82 -151717.2076715877
Lbr82 netRa82 netL82 1.6283385473515223e-10
Rbbr82 netL82 0 320332.57823985495
Cbr82 netL82 0 3.348506201139111e-21

* Branch 83
Rabr83 node_2 netRa83 132180.6654545438
Lbr83 netRa83 netL83 -5.020052708979156e-11
Rbbr83 netL83 0 -160213.71645730478
Cbr83 netL83 0 -2.3699696642370342e-21

* Branch 84
Rabr84 node_2 netRa84 2303802.7231165594
Lbr84 netRa84 netL84 -5.675504131875978e-10
Rbbr84 netL84 0 -2527933.9795251726
Cbr84 netL84 0 -9.743630915490577e-23

* Branch 85
Rabr85 node_2 netRa85 8451084.516057024
Lbr85 netRa85 netL85 -9.418056339807571e-10
Rbbr85 netL85 0 -8630532.16310877
Cbr85 netL85 0 -1.2911525765857581e-23

* Branch 86
Rabr86 node_2 netRa86 -392934.7174822573
Lbr86 netRa86 netL86 2.0672937797386e-10
Rbbr86 netL86 0 495086.1686003746
Cbr86 netL86 0 1.0622735499860059e-21

* Branch 87
Rabr87 node_2 netRa87 839097.8658640755
Lbr87 netRa87 netL87 -3.009194403318253e-10
Rbbr87 netL87 0 -1044894.4764634018
Cbr87 netL87 0 -3.4311584354957066e-22

* Branch 88
Rabr88 node_2 netRa88 107053.14246670993
Lbr88 netRa88 netL88 3.844006312190487e-10
Rbbr88 netL88 0 -2981384.6947413543
Cbr88 netL88 0 1.2081442756622626e-21

* Branch 89
Rabr89 node_2 netRa89 8436.513254550435
Lbr89 netRa89 netL89 -4.0239512169273185e-11
Rbbr89 netL89 0 -631461.8275887589
Cbr89 netL89 0 -7.518195159582029e-21

* Branch 90
Rabr90 node_2 netRa90 542910.6137207444
Lbr90 netRa90 netL90 -2.25014400921659e-10
Rbbr90 netL90 0 -705607.6646728995
Cbr90 netL90 0 -5.871032350303911e-22

* Branch 91
Rabr91 node_2 netRa91 74790.42304794234
Lbr91 netRa91 netL91 4.2294163172695094e-11
Rbbr91 netL91 0 -151631.59274829002
Cbr91 netL91 0 3.732151469495514e-21

* Branch 92
Rabr92 node_2 netRa92 1547686.6360363967
Lbr92 netRa92 netL92 1.0404618396020566e-10
Rbbr92 netL92 0 -1569841.6567262474
Cbr92 netL92 0 4.282988557330728e-23

* Branch 93
Rabr93 node_2 netRa93 397983.90760613297
Lbr93 netRa93 netL93 -2.1240043347360145e-10
Rbbr93 netL93 0 -627897.3223432602
Cbr93 netL93 0 -8.489261323384395e-22

* Branch 94
Rabr94 node_2 netRa94 30473.934785123376
Lbr94 netRa94 netL94 -1.9882243167990436e-11
Rbbr94 netL94 0 -70101.71713706605
Cbr94 netL94 0 -9.292625598189631e-21

* Branch 95
Rabr95 node_2 netRa95 72430.99008863523
Lbr95 netRa95 netL95 -5.488061742896857e-11
Rbbr95 netL95 0 -213749.96799470356
Cbr95 netL95 0 -3.538080163401319e-21

* Branch 96
Rabr96 node_2 netRa96 -7763.718194151846
Lbr96 netRa96 netL96 5.7450719673491367e-11
Rbbr96 netL96 0 388813.0584221618
Cbr96 netL96 0 1.8586086686711387e-20

* Branch 97
Rabr97 node_2 netRa97 -50956.45971217919
Lbr97 netRa97 netL97 -4.4979611008609093e-11
Rbbr97 netL97 0 188482.49807066505
Cbr97 netL97 0 -4.700706058336834e-21

* Branch 98
Rabr98 node_2 netRa98 5461.826638962721
Lbr98 netRa98 netL98 -4.572263280636015e-12
Rbbr98 netL98 0 -7319.35329556302
Cbr98 netL98 0 -1.1390294573504517e-19

* Branch 99
Rabr99 node_2 netRa99 3491818.2500041607
Lbr99 netRa99 netL99 -1.1742032807172028e-10
Rbbr99 netL99 0 -3499001.0135329477
Cbr99 netL99 0 -9.60628313878666e-24

.ends


* Y'23
.subckt yp23 node_2 node_3
* Branch 0
Rabr0 node_2 netRa0 -478.3047431634189
Lbr0 netRa0 netL0 -2.753547515186316e-13
Rbbr0 netL0 node_3 595.8411723412506
Cbr0 netL0 node_3 -9.984478953437894e-19

* Branch 1
Rabr1 node_2 netRa1 -88.5013194496582
Lbr1 netRa1 netL1 1.0783761124904804e-13
Rbbr1 netL1 node_3 229.2778358490099
Cbr1 netL1 node_3 5.051232697940496e-18

* Branch 2
Rabr2 node_2 netRa2 -349.23707594545084
Lbr2 netRa2 netL2 1.5254100562151217e-13
Rbbr2 netL2 node_3 422.4982464524322
Cbr2 netL2 node_3 1.0163204286322895e-18

* Branch 3
Rabr3 node_2 netRa3 -730.5458775817061
Lbr3 netRa3 netL3 2.505285004942009e-13
Rbbr3 netL3 node_3 825.8402629505125
Cbr3 netL3 node_3 4.099868822968035e-19

* Branch 4
Rabr4 node_2 netRa4 -649.6564709275866
Lbr4 netRa4 netL4 5.22376827308577e-13
Rbbr4 netL4 node_3 1110.9315246771134
Cbr4 netL4 node_3 7.030353148743788e-19

* Branch 5
Rabr5 node_2 netRa5 24619.360891874407
Lbr5 netRa5 netL5 6.124728622584321e-12
Rbbr5 netL5 node_3 -28126.33649560077
Cbr5 netL5 node_3 8.909342303960196e-21

* Branch 6
Rabr6 node_2 netRa6 14862.99100181036
Lbr6 netRa6 netL6 -6.2406418729382594e-12
Rbbr6 netL6 node_3 -21245.861405867356
Cbr6 netL6 node_3 -1.9538814632997267e-20

* Branch 7
Rabr7 node_2 netRa7 -217.88525514918146
Lbr7 netRa7 netL7 1.70488394634548e-13
Rbbr7 netL7 node_3 568.6203272829703
Cbr7 netL7 node_3 1.3473554818915548e-18

* Branch 8
Rabr8 node_2 netRa8 24958.27466518607
Lbr8 netRa8 netL8 7.247472652987362e-12
Rbbr8 netL8 node_3 -29961.127931540952
Cbr8 netL8 node_3 9.769224625202167e-21

* Branch 9
Rabr9 node_2 netRa9 -72.48672060840856
Lbr9 netRa9 netL9 1.7374526902251763e-13
Rbbr9 netL9 node_3 1121.5241973878146
Cbr9 netL9 node_3 2.0106448647775515e-18

* Branch 10
Rabr10 node_2 netRa10 53.893488209268845
Lbr10 netRa10 netL10 -1.1330261194755767e-13
Rbbr10 netL10 node_3 -657.5469503927028
Cbr10 netL10 node_3 -3.0375305054412963e-18

* Branch 11
Rabr11 node_2 netRa11 3824.096063352009
Lbr11 netRa11 netL11 -3.335516177662903e-12
Rbbr11 netL11 node_3 -10121.666753867137
Cbr11 netL11 node_3 -8.45240904357392e-20

* Branch 12
Rabr12 node_2 netRa12 1512.9298405895224
Lbr12 netRa12 netL12 -5.326273423325875e-13
Rbbr12 netL12 node_3 -1713.9994217418616
Cbr12 netL12 node_3 -2.0387155942971597e-19

* Branch 13
Rabr13 node_2 netRa13 -23.640550567640368
Lbr13 netRa13 netL13 6.03844963936989e-13
Rbbr13 netL13 node_3 25925.69739492023
Cbr13 netL13 node_3 6.408122855568071e-19

* Branch 14
Rabr14 node_2 netRa14 -17.769607274666285
Lbr14 netRa14 netL14 -1.7148861075222267e-13
Rbbr14 netL14 node_3 3254.8549815512947
Cbr14 netL14 node_3 -3.659434307233372e-18

* Branch 15
Rabr15 node_2 netRa15 -835.0030749380484
Lbr15 netRa15 netL15 9.583764707629898e-13
Rbbr15 netL15 node_3 3768.330491396285
Cbr15 netL15 node_3 2.9787853253970934e-19

* Branch 16
Rabr16 node_2 netRa16 13763.19829718404
Lbr16 netRa16 netL16 5.048786300854284e-12
Rbbr16 netL16 node_3 -17822.66412077138
Cbr16 netL16 node_3 2.072674591356221e-20

* Branch 17
Rabr17 node_2 netRa17 85.89755958757235
Lbr17 netRa17 netL17 -1.3690194012890977e-13
Rbbr17 netL17 node_3 -320.2247852021088
Cbr17 netL17 node_3 -4.836976425509271e-18

* Branch 18
Rabr18 node_2 netRa18 14356.468286071848
Lbr18 netRa18 netL18 -2.5269330274000235e-12
Rbbr18 netL18 node_3 -15517.003129598632
Cbr18 netL18 node_3 -1.13085123778124e-20

* Branch 19
Rabr19 node_2 netRa19 -2688949.8957221946
Lbr19 netRa19 netL19 5.610050015579603e-11
Rbbr19 netL19 node_3 2692550.7146930113
Cbr19 netL19 node_3 7.745775392010991e-24

* Branch 20
Rabr20 node_2 netRa20 1073.6060033325273
Lbr20 netRa20 netL20 5.023555650170802e-13
Rbbr20 netL20 node_3 -1571.1181134217138
Cbr20 netL20 node_3 3.0015921484346553e-19

* Branch 21
Rabr21 node_2 netRa21 1998.2049852904304
Lbr21 netRa21 netL21 5.309494523670794e-12
Rbbr21 netL21 node_3 -37934.453764753984
Cbr21 netL21 node_3 7.327432816799533e-20

* Branch 22
Rabr22 node_2 netRa22 -23.3483691133465
Lbr22 netRa22 netL22 1.6939536666349905e-13
Rbbr22 netL22 node_3 3312.827841670817
Cbr22 netL22 node_3 1.958768982172212e-18

* Branch 23
Rabr23 node_2 netRa23 -2597.3557094541966
Lbr23 netRa23 netL23 3.80902015914156e-12
Rbbr23 netL23 node_3 17770.46695151438
Cbr23 netL23 node_3 8.063086739083614e-20

* Branch 24
Rabr24 node_2 netRa24 137.63894078050666
Lbr24 netRa24 netL24 3.8227851321290454e-13
Rbbr24 netL24 node_3 -3461.56874678711
Cbr24 netL24 node_3 8.38446241145412e-19

* Branch 25
Rabr25 node_2 netRa25 -92508.13060609628
Lbr25 netRa25 netL25 -1.832190737366704e-11
Rbbr25 netL25 node_3 95870.15097445826
Cbr25 netL25 node_3 -2.0722003660208315e-21

* Branch 26
Rabr26 node_2 netRa26 -16.639148064404726
Lbr26 netRa26 netL26 4.0519682057716416e-14
Rbbr26 netL26 node_3 171.00558006579118
Cbr26 netL26 node_3 1.3731688490703913e-17

* Branch 27
Rabr27 node_2 netRa27 -41.48440157830157
Lbr27 netRa27 netL27 1.3968636058126222e-12
Rbbr27 netL27 node_3 42886.33116740388
Cbr27 netL27 node_3 5.196590930350779e-19

* Branch 28
Rabr28 node_2 netRa28 -98.07062933075886
Lbr28 netRa28 netL28 1.9846919542254175e-12
Rbbr28 netL28 node_3 106285.92736927065
Cbr28 netL28 node_3 1.4647973871365833e-19

* Branch 29
Rabr29 node_2 netRa29 -1022.1635760230715
Lbr29 netRa29 netL29 2.5912893269126754e-12
Rbbr29 netL29 node_3 19255.920654050966
Cbr29 netL29 node_3 1.2708033201962625e-19

* Branch 30
Rabr30 node_2 netRa30 -1949.9510227759674
Lbr30 netRa30 netL30 -4.149344830767805e-13
Rbbr30 netL30 node_3 2216.0860590203556
Cbr30 netL30 node_3 -9.629168687232153e-20

* Branch 31
Rabr31 node_2 netRa31 -2875.24871969912
Lbr31 netRa31 netL31 -3.3634971557346723e-12
Rbbr31 netL31 node_3 15469.036163747303
Cbr31 netL31 node_3 -7.680522778577638e-20

* Branch 32
Rabr32 node_2 netRa32 -604.4204987637617
Lbr32 netRa32 netL32 -6.718871241547795e-13
Rbbr32 netL32 node_3 2203.834265083168
Cbr32 netL32 node_3 -5.118300244413803e-19

* Branch 33
Rabr33 node_2 netRa33 -2942.0191747808058
Lbr33 netRa33 netL33 3.5097972315945e-12
Rbbr33 netL33 node_3 7950.448066295672
Cbr33 netL33 node_3 1.4782623065520028e-19

* Branch 34
Rabr34 node_2 netRa34 2872.052047990094
Lbr34 netRa34 netL34 1.2683198077403738e-12
Rbbr34 netL34 node_3 -3849.4244293904276
Cbr34 netL34 node_3 1.1533652558437481e-19

* Branch 35
Rabr35 node_2 netRa35 -28382.768503839015
Lbr35 netRa35 netL35 9.898777815863418e-12
Rbbr35 netL35 node_3 31660.54880228315
Cbr35 netL35 node_3 1.0971873771559593e-20

* Branch 36
Rabr36 node_2 netRa36 -11991551.410429427
Lbr36 netRa36 netL36 2.254704851126276e-10
Rbbr36 netL36 node_3 11995358.328838265
Cbr36 netL36 node_3 1.5671496800501657e-24

* Branch 37
Rabr37 node_2 netRa37 1042.397914623316
Lbr37 netRa37 netL37 -4.1851916149093235e-12
Rbbr37 netL37 node_3 -25847.513887588426
Cbr37 netL37 node_3 -1.4875917490166988e-19

* Branch 38
Rabr38 node_2 netRa38 2263.3116343083134
Lbr38 netRa38 netL38 2.197224633577236e-12
Rbbr38 netL38 node_3 -6476.054476674376
Cbr38 netL38 node_3 1.5145265151872807e-19

* Branch 39
Rabr39 node_2 netRa39 -1477.1256964686863
Lbr39 netRa39 netL39 5.058055509769228e-12
Rbbr39 netL39 node_3 48817.277723373096
Cbr39 netL39 node_3 6.785401801971075e-20

* Branch 40
Rabr40 node_2 netRa40 1402.004721232984
Lbr40 netRa40 netL40 2.353911727707007e-12
Rbbr40 netL40 node_3 -9424.990622587713
Cbr40 netL40 node_3 1.810229539352172e-19

* Branch 41
Rabr41 node_2 netRa41 2233.9808256383694
Lbr41 netRa41 netL41 1.7166263009032465e-12
Rbbr41 netL41 node_3 -4776.755300110823
Cbr41 netL41 node_3 1.6203415433780778e-19

* Branch 42
Rabr42 node_2 netRa42 -8816.571135762382
Lbr42 netRa42 netL42 4.673857063578613e-12
Rbbr42 netL42 node_3 16953.562411614286
Cbr42 netL42 node_3 3.1117037785541566e-20

* Branch 43
Rabr43 node_2 netRa43 -4743.8963805596395
Lbr43 netRa43 netL43 -9.338464222459137e-12
Rbbr43 netL43 node_3 23408.413859157215
Cbr43 netL43 node_3 -8.564682113418493e-20

* Branch 44
Rabr44 node_2 netRa44 0.25557641114557855
Lbr44 netRa44 netL44 -8.887888217478418e-14
Rbbr44 netL44 node_3 -12866.864311340381
Cbr44 netL44 node_3 -6.98214372650022e-18

* Branch 45
Rabr45 node_2 netRa45 2859.812334344375
Lbr45 netRa45 netL45 2.1823420022045407e-12
Rbbr45 netL45 node_3 -5838.199290455357
Cbr45 netL45 node_3 1.31536824163722e-19

* Branch 46
Rabr46 node_2 netRa46 -8176.533503273275
Lbr46 netRa46 netL46 5.6932285546278965e-12
Rbbr46 netL46 node_3 13085.435490965869
Cbr46 netL46 node_3 5.292140014024137e-20

* Branch 47
Rabr47 node_2 netRa47 -5625.748511532648
Lbr47 netRa47 netL47 5.268850194545979e-12
Rbbr47 netL47 node_3 9869.536740477079
Cbr47 netL47 node_3 9.422285712287113e-20

* Branch 48
Rabr48 node_2 netRa48 351.9959317365104
Lbr48 netRa48 netL48 8.742798686814516e-13
Rbbr48 netL48 node_3 -4127.7076482533275
Cbr48 netL48 node_3 6.131434128251345e-19

* Branch 49
Rabr49 node_2 netRa49 -24123.279597530094
Lbr49 netRa49 netL49 7.9753205718513e-12
Rbbr49 netL49 node_3 27718.510120791438
Cbr49 netL49 node_3 1.1899134816045726e-20

* Branch 50
Rabr50 node_2 netRa50 15740.995642051885
Lbr50 netRa50 netL50 6.517026147691974e-12
Rbbr50 netL50 node_3 -18576.982330876577
Cbr50 netL50 node_3 2.2340555428952063e-20

* Branch 51
Rabr51 node_2 netRa51 -22306.090761748175
Lbr51 netRa51 netL51 -3.9843909184385974e-11
Rbbr51 netL51 node_3 194589.8904047049
Cbr51 netL51 node_3 -9.274138358500219e-21

* Branch 52
Rabr52 node_2 netRa52 10026.155756814032
Lbr52 netRa52 netL52 -5.37584737529669e-12
Rbbr52 netL52 node_3 -17443.331228122846
Cbr52 netL52 node_3 -3.06593716137501e-20

* Branch 53
Rabr53 node_2 netRa53 13115.065019818014
Lbr53 netRa53 netL53 6.448673115076745e-12
Rbbr53 netL53 node_3 -18868.644228318757
Cbr53 netL53 node_3 2.6113097930709486e-20

* Branch 54
Rabr54 node_2 netRa54 -123.9246972824507
Lbr54 netRa54 netL54 -1.2801013644312472e-12
Rbbr54 netL54 node_3 20223.703783463006
Cbr54 netL54 node_3 -5.339623446720485e-19

* Branch 55
Rabr55 node_2 netRa55 -19100.432663340744
Lbr55 netRa55 netL55 1.0194891935424332e-11
Rbbr55 netL55 node_3 37296.69699278215
Cbr55 netL55 node_3 1.4280984962884875e-20

* Branch 56
Rabr56 node_2 netRa56 -12286.57458343042
Lbr56 netRa56 netL56 7.847313949161082e-12
Rbbr56 netL56 node_3 18676.575049944982
Cbr56 netL56 node_3 3.41159277535003e-20

* Branch 57
Rabr57 node_2 netRa57 5326.730222315392
Lbr57 netRa57 netL57 9.201205394770424e-12
Rbbr57 netL57 node_3 -21678.57410184309
Cbr57 netL57 node_3 8.018617189065781e-20

* Branch 58
Rabr58 node_2 netRa58 -5541.202091125259
Lbr58 netRa58 netL58 5.56744779031678e-12
Rbbr58 netL58 node_3 12829.144249049625
Cbr58 netL58 node_3 7.805111878404331e-20

* Branch 59
Rabr59 node_2 netRa59 9403.484613096041
Lbr59 netRa59 netL59 -2.3520746432166048e-12
Rbbr59 netL59 node_3 -10381.988703731937
Cbr59 netL59 node_3 -2.4072399597899913e-20

* Branch 60
Rabr60 node_2 netRa60 -1110.6943044979512
Lbr60 netRa60 netL60 5.057662361650065e-12
Rbbr60 netL60 node_3 43205.07571564285
Cbr60 netL60 node_3 1.0406286156804318e-19

* Branch 61
Rabr61 node_2 netRa61 2301.551880120243
Lbr61 netRa61 netL61 6.202802646400402e-12
Rbbr61 netL61 node_3 -36565.53129134542
Cbr61 netL61 node_3 7.420235812245454e-20

* Branch 62
Rabr62 node_2 netRa62 -7546.282377818573
Lbr62 netRa62 netL62 6.897975463228918e-12
Rbbr62 netL62 node_3 15970.004172569354
Cbr62 netL62 node_3 5.710874351213574e-20

* Branch 63
Rabr63 node_2 netRa63 6367.844369104575
Lbr63 netRa63 netL63 4.767461294890257e-12
Rbbr63 netL63 node_3 -13100.711039303495
Cbr63 netL63 node_3 5.724594686742257e-20

* Branch 64
Rabr64 node_2 netRa64 1633.7327228546897
Lbr64 netRa64 netL64 3.3643919123169005e-12
Rbbr64 netL64 node_3 -16044.036181464446
Cbr64 netL64 node_3 1.2890694467688203e-19

* Branch 65
Rabr65 node_2 netRa65 -680537.883317175
Lbr65 netRa65 netL65 -7.215314935174562e-11
Rbbr65 netL65 node_3 698028.8620441228
Cbr65 netL65 node_3 -1.5192297907418301e-22

* Branch 66
Rabr66 node_2 netRa66 649.30003088626
Lbr66 netRa66 netL66 4.595057846687701e-12
Rbbr66 netL66 node_3 -112243.03492486912
Cbr66 netL66 node_3 6.375530482998942e-20

* Branch 67
Rabr67 node_2 netRa67 3579.695397541083
Lbr67 netRa67 netL67 4.588686160306865e-12
Rbbr67 netL67 node_3 -22701.328155696792
Cbr67 netL67 node_3 5.654627698688384e-20

* Branch 68
Rabr68 node_2 netRa68 -4974.039078802437
Lbr68 netRa68 netL68 3.4004145586954565e-12
Rbbr68 netL68 node_3 8410.524978387082
Cbr68 netL68 node_3 8.122880967802767e-20

* Branch 69
Rabr69 node_2 netRa69 -825.4790546788104
Lbr69 netRa69 netL69 1.588830929818913e-12
Rbbr69 netL69 node_3 4326.092063920556
Cbr69 netL69 node_3 4.442123528247369e-19

* Branch 70
Rabr70 node_2 netRa70 -675.8274408185367
Lbr70 netRa70 netL70 1.9051129529947706e-11
Rbbr70 netL70 node_3 211757.58406797657
Cbr70 netL70 node_3 1.3079857884238435e-19

* Branch 71
Rabr71 node_2 netRa71 -655.9899183551734
Lbr71 netRa71 netL71 -8.990256912265097e-13
Rbbr71 netL71 node_3 2669.81448615375
Cbr71 netL71 node_3 -5.136359741439562e-19

* Branch 72
Rabr72 node_2 netRa72 602.7106979269372
Lbr72 netRa72 netL72 1.588464403758068e-11
Rbbr72 netL72 node_3 -177270.44878215567
Cbr72 netL72 node_3 1.5036249344202023e-19

* Branch 73
Rabr73 node_2 netRa73 2247.633515542187
Lbr73 netRa73 netL73 1.2546532902419736e-11
Rbbr73 netL73 node_3 -32776.77826487445
Cbr73 netL73 node_3 1.7065477748592993e-19

* Branch 74
Rabr74 node_2 netRa74 2800.628172933735
Lbr74 netRa74 netL74 1.0459325093790525e-11
Rbbr74 netL74 node_3 -20515.420319740315
Cbr74 netL74 node_3 1.821916069585832e-19

* Branch 75
Rabr75 node_2 netRa75 1805.11097274485
Lbr75 netRa75 netL75 4.288585719604714e-12
Rbbr75 netL75 node_3 -10302.261496416913
Cbr75 netL75 node_3 2.3063142667524927e-19

* Branch 76
Rabr76 node_2 netRa76 -3593.873826193797
Lbr76 netRa76 netL76 1.000704947160422e-11
Rbbr76 netL76 node_3 16727.407298278962
Cbr76 netL76 node_3 1.66433654325129e-19

* Branch 77
Rabr77 node_2 netRa77 3180.8547260289197
Lbr77 netRa77 netL77 5.048215879801241e-12
Rbbr77 netL77 node_3 -9496.866290888822
Cbr77 netL77 node_3 1.671364754598797e-19

* Branch 78
Rabr78 node_2 netRa78 1174.633032797861
Lbr78 netRa78 netL78 4.882495723677448e-12
Rbbr78 netL78 node_3 -16718.17917547651
Cbr78 netL78 node_3 2.489295311245841e-19

* Branch 79
Rabr79 node_2 netRa79 -112335.01478382996
Lbr79 netRa79 netL79 -3.7143579482325046e-11
Rbbr79 netL79 node_3 118354.33923447409
Cbr79 netL79 node_3 -2.794026490879308e-21

* Branch 80
Rabr80 node_2 netRa80 -585.6231271699074
Lbr80 netRa80 netL80 1.5334752827581992e-12
Rbbr80 netL80 node_3 6445.711657420153
Cbr80 netL80 node_3 4.058925690189842e-19

* Branch 81
Rabr81 node_2 netRa81 -7182.320132880563
Lbr81 netRa81 netL81 -1.0564197173264506e-11
Rbbr81 netL81 node_3 15098.755237228435
Cbr81 netL81 node_3 -9.747633346738067e-20

* Branch 82
Rabr82 node_2 netRa82 -1418.6930475274548
Lbr82 netRa82 netL82 -7.189292975159398e-12
Rbbr82 netL82 node_3 20723.663300408654
Cbr82 netL82 node_3 -2.4510793211886996e-19

* Branch 83
Rabr83 node_2 netRa83 -1648.7112869888117
Lbr83 netRa83 netL83 -6.928040421241032e-12
Rbbr83 netL83 node_3 17654.26470460187
Cbr83 netL83 node_3 -2.3862602642693787e-19

* Branch 84
Rabr84 node_2 netRa84 -801.091472484966
Lbr84 netRa84 netL84 -5.602601584127297e-12
Rbbr84 netL84 node_3 27359.90744826456
Cbr84 netL84 node_3 -2.5686072058676374e-19

* Branch 85
Rabr85 node_2 netRa85 -650.5208823131106
Lbr85 netRa85 netL85 -5.404050459810162e-12
Rbbr85 netL85 node_3 30127.92883637768
Cbr85 netL85 node_3 -2.774179908750616e-19

* Branch 86
Rabr86 node_2 netRa86 -4167.671617214262
Lbr86 netRa86 netL86 -8.286477497149431e-12
Rbbr86 netL86 node_3 15663.202506132395
Cbr86 netL86 node_3 -1.2712773648722517e-19

* Branch 87
Rabr87 node_2 netRa87 -2333.120141408307
Lbr87 netRa87 netL87 -6.987972869080174e-12
Rbbr87 netL87 node_3 14258.632502454479
Cbr87 netL87 node_3 -2.105395960431139e-19

* Branch 88
Rabr88 node_2 netRa88 -770.8314132032795
Lbr88 netRa88 netL88 -5.518502986367294e-12
Rbbr88 netL88 node_3 25844.425551201613
Cbr88 netL88 node_3 -2.7858316616763667e-19

* Branch 89
Rabr89 node_2 netRa89 -1244.1603951521813
Lbr89 netRa89 netL89 -5.923969010252754e-12
Rbbr89 netL89 node_3 18512.738808100825
Cbr89 netL89 node_3 -2.582014691994357e-19

* Branch 90
Rabr90 node_2 netRa90 -2076.381770483417
Lbr90 netRa90 netL90 -6.598148463852055e-12
Rbbr90 netL90 node_3 14457.603846338148
Cbr90 netL90 node_3 -2.203742506811265e-19

* Branch 91
Rabr91 node_2 netRa91 -4512.276153870292
Lbr91 netRa91 netL91 8.697166292785183e-12
Rbbr91 netL91 node_3 16925.807138400225
Cbr91 netL91 node_3 1.136808275080501e-19

* Branch 92
Rabr92 node_2 netRa92 -394242.31061088765
Lbr92 netRa92 netL92 -8.088906342174706e-11
Rbbr92 netL92 node_3 406178.7965594013
Cbr92 netL92 node_3 -5.052343408406476e-22

* Branch 93
Rabr93 node_2 netRa93 167.90304286175905
Lbr93 netRa93 netL93 3.5247785057610793e-12
Rbbr93 netL93 node_3 -61562.37377273505
Cbr93 netL93 node_3 3.48828900441195e-19

* Branch 94
Rabr94 node_2 netRa94 -18182.373705873357
Lbr94 netRa94 netL94 -5.267875213776276e-12
Rbbr94 netL94 node_3 23036.538148196323
Cbr94 netL94 node_3 -1.258318999714772e-20

* Branch 95
Rabr95 node_2 netRa95 -667.9465495002913
Lbr95 netRa95 netL95 5.650735209364596e-12
Rbbr95 netL95 node_3 151550.56615640697
Cbr95 netL95 node_3 5.49709350910869e-20

* Branch 96
Rabr96 node_2 netRa96 -202405.49481672095
Lbr96 netRa96 netL96 1.3639261452698855e-11
Rbbr96 netL96 node_3 205712.2018151857
Cbr96 netL96 node_3 3.274377677083449e-22

* Branch 97
Rabr97 node_2 netRa97 313.32450779213093
Lbr97 netRa97 netL97 -1.6032612735759053e-13
Rbbr97 netL97 node_3 -557.7247347558888
Cbr97 netL97 node_3 -9.12035672533221e-19

* Branch 98
Rabr98 node_2 netRa98 145.15809502739847
Lbr98 netRa98 netL98 -1.9701370991769804e-13
Rbbr98 netL98 node_3 -843.0360523423915
Cbr98 netL98 node_3 -1.557126623081833e-18

* Branch 99
Rabr99 node_2 netRa99 171.68638190998706
Lbr99 netRa99 netL99 -9.617070708865369e-14
Rbbr99 netL99 node_3 -231.96318368267262
Cbr99 netL99 node_3 -2.374268159834037e-18

.ends


* Y'24
.subckt yp24 node_2 node_4
* Branch 0
Rabr0 node_2 netRa0 -40.69069699598561
Lbr0 netRa0 netL0 -3.053494933553719e-14
Rbbr0 netL0 node_4 67.83645780858558
Cbr0 netL0 node_4 -1.154256057718543e-17

* Branch 1
Rabr1 node_2 netRa1 13.792912690545185
Lbr1 netRa1 netL1 4.0498469297802516e-14
Rbbr1 netL1 node_4 -109.39730827588181
Cbr1 netL1 node_4 3.1787112833334116e-17

* Branch 2
Rabr2 node_2 netRa2 8856.537575877674
Lbr2 netRa2 netL2 -7.22586672649553e-13
Rbbr2 netL2 node_4 -8923.052466472955
Cbr2 netL2 node_4 -9.104145899198707e-21

* Branch 3
Rabr3 node_2 netRa3 757.9322493270797
Lbr3 netRa3 netL3 -9.067786274843665e-14
Rbbr3 netL3 node_4 -770.1105220260981
Cbr3 netL3 node_4 -1.5439676098933712e-19

* Branch 4
Rabr4 node_2 netRa4 2.586020554074472
Lbr4 netRa4 netL4 6.917383489514438e-15
Rbbr4 netL4 node_4 -26.572376436005165
Cbr4 netL4 node_4 1.150053534326043e-16

* Branch 5
Rabr5 node_2 netRa5 -53.403670945541094
Lbr5 netRa5 netL5 -3.5446025397722146e-12
Rbbr5 netL5 node_4 -913267.7727005405
Cbr5 netL5 node_4 -8.486442432706384e-20

* Branch 6
Rabr6 node_2 netRa6 -2717.3699356808143
Lbr6 netRa6 netL6 -3.20296061483672e-13
Rbbr6 netL6 node_4 2734.6260750818656
Cbr6 netL6 node_4 -4.3241994731068426e-20

* Branch 7
Rabr7 node_2 netRa7 4130.100684027088
Lbr7 netRa7 netL7 1.1567332762779524e-12
Rbbr7 netL7 node_4 -4906.99767521015
Cbr7 netL7 node_4 5.75064123966168e-20

* Branch 8
Rabr8 node_2 netRa8 -11.101801206634683
Lbr8 netRa8 netL8 -5.794985409491733e-14
Rbbr8 netL8 node_4 411.1479367883547
Cbr8 netL8 node_4 -1.469397491139398e-17

* Branch 9
Rabr9 node_2 netRa9 -48.567073204606274
Lbr9 netRa9 netL9 6.850921080437741e-14
Rbbr9 netL9 node_4 151.20657417731113
Cbr9 netL9 node_4 9.002196621033316e-18

* Branch 10
Rabr10 node_2 netRa10 -705.4297407858113
Lbr10 netRa10 netL10 -3.718305041227725e-13
Rbbr10 netL10 node_4 1265.592055035245
Cbr10 netL10 node_4 -4.217001511716304e-19

* Branch 11
Rabr11 node_2 netRa11 -18690.679104133535
Lbr11 netRa11 netL11 1.3328939846332905e-12
Rbbr11 netL11 node_4 18950.487619748947
Cbr11 netL11 node_4 3.757058928873324e-21

* Branch 12
Rabr12 node_2 netRa12 119.48143643056486
Lbr12 netRa12 netL12 5.588475303139147e-14
Rbbr12 netL12 node_4 -189.16282696937898
Cbr12 netL12 node_4 2.499080563580573e-18

* Branch 13
Rabr13 node_2 netRa13 -36866.15587786138
Lbr13 netRa13 netL13 2.158978066169015e-12
Rbbr13 netL13 node_4 37002.05773274887
Cbr13 netL13 node_4 1.5806156891138387e-21

* Branch 14
Rabr14 node_2 netRa14 17523.811714202846
Lbr14 netRa14 netL14 6.06921605737336e-12
Rbbr14 netL14 node_4 -19555.711204013573
Cbr14 netL14 node_4 1.784441612328526e-20

* Branch 15
Rabr15 node_2 netRa15 3273.751783691772
Lbr15 netRa15 netL15 2.423834612499989e-12
Rbbr15 netL15 node_4 -7492.892590237229
Cbr15 netL15 node_4 1.0038024460886354e-19

* Branch 16
Rabr16 node_2 netRa16 -271805.09719859954
Lbr16 netRa16 netL16 -2.6479023881601953e-11
Rbbr16 netL16 node_4 277581.3184353983
Cbr16 netL16 node_4 -3.5159232912382446e-22

* Branch 17
Rabr17 node_2 netRa17 874.2488928636468
Lbr17 netRa17 netL17 1.0609049529976941e-12
Rbbr17 netL17 node_4 -4177.397166712725
Cbr17 netL17 node_4 2.9705848320378636e-19

* Branch 18
Rabr18 node_2 netRa18 44.67517157607244
Lbr18 netRa18 netL18 2.4199016027509468e-14
Rbbr18 netL18 node_4 -71.5365686707761
Cbr18 netL18 node_4 7.646618984071468e-18

* Branch 19
Rabr19 node_2 netRa19 28.192601040809443
Lbr19 netRa19 netL19 1.151109303477133e-13
Rbbr19 netL19 node_4 -1033.1918890186334
Cbr19 netL19 node_4 4.260434535706262e-18

* Branch 20
Rabr20 node_2 netRa20 -72.26552760424875
Lbr20 netRa20 netL20 2.006926928291624e-13
Rbbr20 netL20 node_4 1450.0477586848058
Cbr20 netL20 node_4 1.826591869993526e-18

* Branch 21
Rabr21 node_2 netRa21 -25.510695368599713
Lbr21 netRa21 netL21 -1.715733090598778e-14
Rbbr21 netL21 node_4 56.81272109759397
Cbr21 netL21 node_4 -1.1977871505832493e-17

* Branch 22
Rabr22 node_2 netRa22 151.23575174197182
Lbr22 netRa22 netL22 3.251810772066715e-13
Rbbr22 netL22 node_4 -1556.0325796961038
Cbr22 netL22 node_4 1.4343504334974922e-18

* Branch 23
Rabr23 node_2 netRa23 -348292.65637846896
Lbr23 netRa23 netL23 -1.1356803053704135e-11
Rbbr23 netL23 node_4 349089.1316378933
Cbr23 netL23 node_4 -9.34572497517335e-23

* Branch 24
Rabr24 node_2 netRa24 13.785301123485658
Lbr24 netRa24 netL24 -1.9522887581951457e-13
Rbbr24 netL24 node_4 -3478.234212602736
Cbr24 netL24 node_4 -3.2915575855042262e-18

* Branch 25
Rabr25 node_2 netRa25 3266.516814435491
Lbr25 netRa25 netL25 -1.8253252470949037e-12
Rbbr25 netL25 node_4 -5723.610269081174
Cbr25 netL25 node_4 -9.67576764999674e-20

* Branch 26
Rabr26 node_2 netRa26 625590.4504771926
Lbr26 netRa26 netL26 1.1823242874666875e-11
Rbbr26 netL26 node_4 -625962.7549209903
Cbr26 netL26 node_4 3.020139642178992e-23

* Branch 27
Rabr27 node_2 netRa27 -3989.1294207907713
Lbr27 netRa27 netL27 -4.869725793691067e-13
Rbbr27 netL27 node_4 4082.8660171118986
Cbr27 netL27 node_4 -2.9956376824838075e-20

* Branch 28
Rabr28 node_2 netRa28 -9.20096486967337
Lbr28 netRa28 netL28 -1.3042035356344887e-14
Rbbr28 netL28 node_4 47.88268219819259
Cbr28 netL28 node_4 -3.026820986820458e-17

* Branch 29
Rabr29 node_2 netRa29 -7.465378229808578
Lbr29 netRa29 netL29 1.4008265589976557e-14
Rbbr29 netL29 node_4 18.75510579725338
Cbr29 netL29 node_4 9.723806620389398e-17

* Branch 30
Rabr30 node_2 netRa30 -698.018196966947
Lbr30 netRa30 netL30 -3.8987552076530413e-13
Rbbr30 netL30 node_4 1362.1779720737607
Cbr30 netL30 node_4 -4.1357895979368805e-19

* Branch 31
Rabr31 node_2 netRa31 -129.68180142236136
Lbr31 netRa31 netL31 9.394122766487039e-13
Rbbr31 netL31 node_4 7533.390424860997
Cbr31 netL31 node_4 8.674061173405387e-19

* Branch 32
Rabr32 node_2 netRa32 929.6222502107798
Lbr32 netRa32 netL32 -1.083387026248589e-12
Rbbr32 netL32 node_4 -2027.716822571995
Cbr32 netL32 node_4 -5.6514324390241745e-19

* Branch 33
Rabr33 node_2 netRa33 86618.0782704315
Lbr33 netRa33 netL33 -1.4285668937286811e-11
Rbbr33 netL33 node_4 -94211.5549058533
Cbr33 netL33 node_4 -1.7464929508359835e-21

* Branch 34
Rabr34 node_2 netRa34 79.01547007546375
Lbr34 netRa34 netL34 4.552834153077596e-13
Rbbr34 netL34 node_4 -5010.372813096916
Cbr34 netL34 node_4 1.253001197518132e-18

* Branch 35
Rabr35 node_2 netRa35 -44.24050054681007
Lbr35 netRa35 netL35 -2.3181635865383613e-12
Rbbr35 netL35 node_4 1533817.523544897
Cbr35 netL35 node_4 -1.2568901635981568e-19

* Branch 36
Rabr36 node_2 netRa36 24.019551581994364
Lbr36 netRa36 netL36 5.5116048871356244e-14
Rbbr36 netL36 node_4 -258.47665766496215
Cbr36 netL36 node_4 9.161256580377683e-18

* Branch 37
Rabr37 node_2 netRa37 44.550119895413395
Lbr37 netRa37 netL37 5.109205123026833e-14
Rbbr37 netL37 node_4 -232.39446341733907
Cbr37 netL37 node_4 5.010334075744296e-18

* Branch 38
Rabr38 node_2 netRa38 -1131.5932150796475
Lbr38 netRa38 netL38 1.1237648330686458e-12
Rbbr38 netL38 node_4 2501.9725369384787
Cbr38 netL38 node_4 3.9202191238503473e-19

* Branch 39
Rabr39 node_2 netRa39 1617.6415107588953
Lbr39 netRa39 netL39 3.406821368837283e-13
Rbbr39 netL39 node_4 -1845.921821408865
Cbr39 netL39 node_4 1.1438728257600054e-19

* Branch 40
Rabr40 node_2 netRa40 5.22738700541949
Lbr40 netRa40 netL40 2.199191962335892e-14
Rbbr40 netL40 node_4 -162.26382657958004
Cbr40 netL40 node_4 2.7309146407963883e-17

* Branch 41
Rabr41 node_2 netRa41 -2193.9210613027813
Lbr41 netRa41 netL41 3.4834562789259967e-12
Rbbr41 netL41 node_4 17825.76332014207
Cbr41 netL41 node_4 8.746632499878494e-20

* Branch 42
Rabr42 node_2 netRa42 -311.19294985784364
Lbr42 netRa42 netL42 2.661012037465977e-13
Rbbr42 netL42 node_4 604.2488205307384
Cbr42 netL42 node_4 1.4018489984151556e-18

* Branch 43
Rabr43 node_2 netRa43 121.19713630427572
Lbr43 netRa43 netL43 2.058707927720395e-13
Rbbr43 netL43 node_4 -590.7871291712383
Cbr43 netL43 node_4 2.9252103938620943e-18

* Branch 44
Rabr44 node_2 netRa44 -812.0107054727043
Lbr44 netRa44 netL44 1.159314544755144e-12
Rbbr44 netL44 node_4 5448.430989030857
Cbr44 netL44 node_4 2.5839568787892464e-19

* Branch 45
Rabr45 node_2 netRa45 -15354.27316068673
Lbr45 netRa45 netL45 -8.121550329265582e-12
Rbbr45 netL45 node_4 24845.119082938916
Cbr45 netL45 node_4 -2.1394057794031156e-20

* Branch 46
Rabr46 node_2 netRa46 149.97195382105556
Lbr46 netRa46 netL46 3.5501682639922534e-14
Rbbr46 netL46 node_4 -172.50523518189922
Cbr46 netL46 node_4 1.3752088291364175e-18

* Branch 47
Rabr47 node_2 netRa47 2593421.532200781
Lbr47 netRa47 netL47 3.9177176296280365e-11
Rbbr47 netL47 node_4 -2595187.88111517
Cbr47 netL47 node_4 5.821706785204226e-24

* Branch 48
Rabr48 node_2 netRa48 887439.1672571623
Lbr48 netRa48 netL48 -2.809784767861319e-11
Rbbr48 netL48 node_4 -888658.9390124234
Cbr48 netL48 node_4 -3.561865184375347e-23

* Branch 49
Rabr49 node_2 netRa49 52.14159950459864
Lbr49 netRa49 netL49 -1.0315173614836706e-13
Rbbr49 netL49 node_4 -414.52955014226757
Cbr49 netL49 node_4 -4.690462774921806e-18

* Branch 50
Rabr50 node_2 netRa50 -220445.86564350565
Lbr50 netRa50 netL50 -1.518604978229901e-11
Rbbr50 netL50 node_4 221539.1236553219
Cbr50 netL50 node_4 -3.111342990571496e-22

* Branch 51
Rabr51 node_2 netRa51 11752.329674275074
Lbr51 netRa51 netL51 4.939665680948187e-12
Rbbr51 netL51 node_4 -13559.744665915441
Cbr51 netL51 node_4 3.110672520748591e-20

* Branch 52
Rabr52 node_2 netRa52 10491.134009001273
Lbr52 netRa52 netL52 8.171622545239358e-12
Rbbr52 netL52 node_4 -32115.82422665691
Cbr52 netL52 node_4 2.4401785731482072e-20

* Branch 53
Rabr53 node_2 netRa53 -1145.8341741154577
Lbr53 netRa53 netL53 2.175730729602082e-12
Rbbr53 netL53 node_4 13623.396372106796
Cbr53 netL53 node_4 1.373883582221923e-19

* Branch 54
Rabr54 node_2 netRa54 2.9625313917285183
Lbr54 netRa54 netL54 -4.6246001623442276e-14
Rbbr54 netL54 node_4 -1054.779767797064
Cbr54 netL54 node_4 -1.330576699741414e-17

* Branch 55
Rabr55 node_2 netRa55 -1324.572546468359
Lbr55 netRa55 netL55 1.960318899886046e-12
Rbbr55 netL55 node_4 5426.591730706051
Cbr55 netL55 node_4 2.70120551983308e-19

* Branch 56
Rabr56 node_2 netRa56 -542.9373065693563
Lbr56 netRa56 netL56 5.076069934001196e-13
Rbbr56 netL56 node_4 1376.526519017477
Cbr56 netL56 node_4 6.751394899523644e-19

* Branch 57
Rabr57 node_2 netRa57 -312910.5267029986
Lbr57 netRa57 netL57 -1.5920528828349502e-11
Rbbr57 netL57 node_4 313945.10830319
Cbr57 netL57 node_4 -1.6211447697991097e-22

* Branch 58
Rabr58 node_2 netRa58 450.0776938829696
Lbr58 netRa58 netL58 -5.796112536808805e-13
Rbbr58 netL58 node_4 -1815.2103119444237
Cbr58 netL58 node_4 -7.042690756568516e-19

* Branch 59
Rabr59 node_2 netRa59 -1293.1882120094838
Lbr59 netRa59 netL59 8.108539481146203e-13
Rbbr59 netL59 node_4 2361.6349863142163
Cbr59 netL59 node_4 2.6462970551620745e-19

* Branch 60
Rabr60 node_2 netRa60 1166336.331003357
Lbr60 netRa60 netL60 -4.0850890719357385e-10
Rbbr60 netL60 node_4 -1309113.5087804561
Cbr60 netL60 node_4 -2.6707612101292753e-22

* Branch 61
Rabr61 node_2 netRa61 27685.911178483868
Lbr61 netRa61 netL61 -6.117147688624099e-12
Rbbr61 netL61 node_4 -30229.498112343204
Cbr61 netL61 node_4 -7.301479898532184e-21

* Branch 62
Rabr62 node_2 netRa62 13105.497587182064
Lbr62 netRa62 netL62 3.2392398311428162e-12
Rbbr62 netL62 node_4 -14181.508054367503
Cbr62 netL62 node_4 1.7446812862585004e-20

* Branch 63
Rabr63 node_2 netRa63 244.1218550341246
Lbr63 netRa63 netL63 -1.013604102413227e-12
Rbbr63 netL63 node_4 -3678.237793424686
Cbr63 netL63 node_4 -1.1109674144866299e-18

* Branch 64
Rabr64 node_2 netRa64 -2913.847477297522
Lbr64 netRa64 netL64 -4.386698326374838e-12
Rbbr64 netL64 node_4 8881.01523785176
Cbr64 netL64 node_4 -1.704438464169224e-19

* Branch 65
Rabr65 node_2 netRa65 -17427.63565859852
Lbr65 netRa65 netL65 -1.1614011683625884e-11
Rbbr65 netL65 node_4 25334.36974681018
Cbr65 netL65 node_4 -2.6351767908393572e-20

* Branch 66
Rabr66 node_2 netRa66 32.8196323550093
Lbr66 netRa66 netL66 1.3732506145919187e-12
Rbbr66 netL66 node_4 -92736.71772906417
Cbr66 netL66 node_4 5.011559209655011e-19

* Branch 67
Rabr67 node_2 netRa67 -4174.890240650708
Lbr67 netRa67 netL67 -9.263547822429073e-13
Rbbr67 netL67 node_4 4503.906329419793
Cbr67 netL67 node_4 -4.929125817179781e-20

* Branch 68
Rabr68 node_2 netRa68 -5835.406027913423
Lbr68 netRa68 netL68 -6.939350701960113e-12
Rbbr68 netL68 node_4 25580.888428738428
Cbr68 netL68 node_4 -4.661096105831774e-20

* Branch 69
Rabr69 node_2 netRa69 -285.158442197059
Lbr69 netRa69 netL69 2.636553613155615e-12
Rbbr69 netL69 node_4 61500.14118184535
Cbr69 netL69 node_4 1.4809275983123889e-19

* Branch 70
Rabr70 node_2 netRa70 34.466059609378284
Lbr70 netRa70 netL70 9.987459221292848e-14
Rbbr70 netL70 node_4 -628.517494006292
Cbr70 netL70 node_4 4.63069671757077e-18

* Branch 71
Rabr71 node_2 netRa71 -114.79519780699927
Lbr71 netRa71 netL71 6.571641513787072e-13
Rbbr71 netL71 node_4 7855.485291869779
Cbr71 netL71 node_4 7.227668569945987e-19

* Branch 72
Rabr72 node_2 netRa72 20040.74710971411
Lbr72 netRa72 netL72 -1.5955669116123123e-10
Rbbr72 netL72 node_4 -2907799.3607186116
Cbr72 netL72 node_4 -2.7118006820252963e-21

* Branch 73
Rabr73 node_2 netRa73 171.69379067877475
Lbr73 netRa73 netL73 -1.4906805108242643e-12
Rbbr73 netL73 node_4 -10274.168482096522
Cbr73 netL73 node_4 -8.373553390489603e-19

* Branch 74
Rabr74 node_2 netRa74 -16.105959249099413
Lbr74 netRa74 netL74 -1.7964448833813425e-12
Rbbr74 netL74 node_4 160754.74824473338
Cbr74 netL74 node_4 -7.279391040196011e-19

* Branch 75
Rabr75 node_2 netRa75 -1678.5217043670093
Lbr75 netRa75 netL75 6.257719603001073e-12
Rbbr75 netL75 node_4 13997.0545461165
Cbr75 netL75 node_4 2.659787499030441e-19

* Branch 76
Rabr76 node_2 netRa76 -1865.6566664288268
Lbr76 netRa76 netL76 4.83131761136026e-12
Rbbr76 netL76 node_4 8234.653873159572
Cbr76 netL76 node_4 3.14192138484606e-19

* Branch 77
Rabr77 node_2 netRa77 -1178.6773893225543
Lbr77 netRa77 netL77 1.0635239615508365e-11
Rbbr77 netL77 node_4 53664.293574700234
Cbr77 netL77 node_4 1.6768758273492467e-19

* Branch 78
Rabr78 node_2 netRa78 -6253.754061325107
Lbr78 netRa78 netL78 1.518695023181843e-12
Rbbr78 netL78 node_4 6420.190086020494
Cbr78 netL78 node_4 3.782256219584885e-20

* Branch 79
Rabr79 node_2 netRa79 -1291.8404935622457
Lbr79 netRa79 netL79 3.851375357419464e-12
Rbbr79 netL79 node_4 18222.387874161155
Cbr79 netL79 node_4 1.6347476042643355e-19

* Branch 80
Rabr80 node_2 netRa80 -12193.018298515117
Lbr80 netRa80 netL80 -2.5438978596468853e-12
Rbbr80 netL80 node_4 13858.134966683545
Cbr80 netL80 node_4 -1.505589613741325e-20

* Branch 81
Rabr81 node_2 netRa81 8110.871600307694
Lbr81 netRa81 netL81 1.8763697679437486e-11
Rbbr81 netL81 node_4 -32794.14158070497
Cbr81 netL81 node_4 7.057487402361208e-20

* Branch 82
Rabr82 node_2 netRa82 -2.299266309455947
Lbr82 netRa82 netL82 -1.1405073898560635e-12
Rbbr82 netL82 node_4 484536.562790308
Cbr82 netL82 node_4 -1.0827879895139395e-18

* Branch 83
Rabr83 node_2 netRa83 -2151.8618042039843
Lbr83 netRa83 netL83 3.8335966575469154e-12
Rbbr83 netL83 node_4 5502.178917283708
Cbr83 netL83 node_4 3.237237912560736e-19

* Branch 84
Rabr84 node_2 netRa84 33856.25019709521
Lbr84 netRa84 netL84 2.6547196072408177e-11
Rbbr84 netL84 node_4 -46111.905924744344
Cbr84 netL84 node_4 1.7005304396877514e-20

* Branch 85
Rabr85 node_2 netRa85 5196.12979249994
Lbr85 netRa85 netL85 1.268956463480302e-11
Rbbr85 netL85 node_4 -24093.43858094189
Cbr85 netL85 node_4 1.0140170609500975e-19

* Branch 86
Rabr86 node_2 netRa86 -197.2344477314641
Lbr86 netRa86 netL86 -1.8800967479569113e-12
Rbbr86 netL86 node_4 13512.26453406436
Cbr86 netL86 node_4 -7.070936699262517e-19

* Branch 87
Rabr87 node_2 netRa87 708.9953323972161
Lbr87 netRa87 netL87 4.9132336706539145e-12
Rbbr87 netL87 node_4 -103684.25995131441
Cbr87 netL87 node_4 6.69617442947027e-20

* Branch 88
Rabr88 node_2 netRa88 -1769.7099993768045
Lbr88 netRa88 netL88 9.244749204917251e-12
Rbbr88 netL88 node_4 32173.10899519209
Cbr88 netL88 node_4 1.620586094797055e-19

* Branch 89
Rabr89 node_2 netRa89 -213.70484638690615
Lbr89 netRa89 netL89 -2.193472129013422e-12
Rbbr89 netL89 node_4 16464.818142660588
Cbr89 netL89 node_4 -6.262588804302396e-19

* Branch 90
Rabr90 node_2 netRa90 -16869.971741165784
Lbr90 netRa90 netL90 1.5017560117143312e-11
Rbbr90 netL90 node_4 25586.676559984124
Cbr90 netL90 node_4 3.4776447665779376e-20

* Branch 91
Rabr91 node_2 netRa91 -514.7320063953274
Lbr91 netRa91 netL91 -3.784515283177251e-12
Rbbr91 netL91 node_4 19957.53734844837
Cbr91 netL91 node_4 -3.697123783072095e-19

* Branch 92
Rabr92 node_2 netRa92 2845.5510899995525
Lbr92 netRa92 netL92 2.8698654530962166e-12
Rbbr92 netL92 node_4 -4211.490751462103
Cbr92 netL92 node_4 2.3959440459347452e-19

* Branch 93
Rabr93 node_2 netRa93 -15841.272823039038
Lbr93 netRa93 netL93 -1.4312047143929091e-11
Rbbr93 netL93 node_4 24562.89915869587
Cbr93 netL93 node_4 -3.679900944898913e-20

* Branch 94
Rabr94 node_2 netRa94 -1539.0823208667805
Lbr94 netRa94 netL94 -9.905939864517732e-12
Rbbr94 netL94 node_4 218902.50628612135
Cbr94 netL94 node_4 -2.950404930204975e-20

* Branch 95
Rabr95 node_2 netRa95 -701.3455833688738
Lbr95 netRa95 netL95 -1.3079309440030155e-13
Rbbr95 netL95 node_4 766.6159108574544
Cbr95 netL95 node_4 -2.4341709576175307e-19

* Branch 96
Rabr96 node_2 netRa96 117529.01607311184
Lbr96 netRa96 netL96 -7.227656963856597e-12
Rbbr96 netL96 node_4 -119136.86515917444
Cbr96 netL96 node_4 -5.158721900586212e-22

* Branch 97
Rabr97 node_2 netRa97 12.688566054267984
Lbr97 netRa97 netL97 -1.4303905207869374e-14
Rbbr97 netL97 node_4 -19.730647559888027
Cbr97 netL97 node_4 -5.621675401896894e-17

* Branch 98
Rabr98 node_2 netRa98 -58.61641436419651
Lbr98 netRa98 netL98 -4.302831076536464e-14
Rbbr98 netL98 node_4 159.6918062869338
Cbr98 netL98 node_4 -4.651834024039142e-18

* Branch 99
Rabr99 node_2 netRa99 -8.26726060668454
Lbr99 netRa99 netL99 -9.107189806760893e-15
Rbbr99 netL99 node_4 20.48656631702315
Cbr99 netL99 node_4 -5.75874690158364e-17

.ends


* Y'33
.subckt yp33 node_3 0
* Branch 0
Rabr0 node_3 netRa0 0.31961066117420983
Lbr0 netRa0 netL0 -2.1655922281829162e-16
Rbbr0 netL0 0 -0.3989136745100733
Cbr0 netL0 0 -1.605947119829523e-15

* Branch 1
Rabr1 node_3 netRa1 0.14358174638989338
Lbr1 netRa1 netL1 -2.705090749965482e-16
Rbbr1 netL1 0 -0.397520654886607
Cbr1 netL1 0 -4.1050257883092245e-15

* Branch 2
Rabr2 node_3 netRa2 -0.8049686151148164
Lbr2 netRa2 netL2 3.4302866736168657e-16
Rbbr2 netL2 0 0.8851278514095338
Cbr2 netL2 0 4.661556900692231e-16

* Branch 3
Rabr3 node_3 netRa3 -0.06546017364404173
Lbr3 netRa3 netL3 -1.300590893033745e-15
Rbbr3 netL3 0 -33.79270606184586
Cbr3 netL3 0 -1.4263016819811441e-15

* Branch 4
Rabr4 node_3 netRa4 0.041831190995913196
Lbr4 netRa4 netL4 -1.0942706335048059e-16
Rbbr4 netL4 0 -0.1997758833627107
Cbr4 netL4 0 -1.1046399814656894e-14

* Branch 5
Rabr5 node_3 netRa5 -1.14603920417318
Lbr5 netRa5 netL5 -2.882919409421292e-16
Rbbr5 netL5 0 1.194215629491266
Cbr5 netL5 0 -2.1432001020956252e-16

* Branch 6
Rabr6 node_3 netRa6 256.2121590407966
Lbr6 netRa6 netL6 7.182291485212335e-15
Rbbr6 netL6 0 -256.3437005536806
Cbr6 netL6 0 1.0953575868485987e-19

* Branch 7
Rabr7 node_3 netRa7 -15.822553082397093
Lbr7 netRa7 netL7 6.021871914196894e-15
Rbbr7 netL7 0 17.14109932801034
Cbr7 netL7 0 2.1733870845194877e-17

* Branch 8
Rabr8 node_3 netRa8 -1159.6731533316329
Lbr8 netRa8 netL8 -5.793480967132485e-13
Rbbr8 netL8 0 1441.2580176225824
Cbr8 netL8 0 -3.555144834183334e-19

* Branch 9
Rabr9 node_3 netRa9 -26948.74056126224
Lbr9 netRa9 netL9 1.1648788679853134e-11
Rbbr9 netL9 0 28906.7764130406
Cbr9 netL9 0 1.466807548298971e-20

* Branch 10
Rabr10 node_3 netRa10 403.6316901675677
Lbr10 netRa10 netL10 -3.207670890245981e-13
Rbbr10 netL10 0 -519.0950445898014
Cbr10 netL10 0 -1.4805090141297743e-18

* Branch 11
Rabr11 node_3 netRa11 -78.61808803936636
Lbr11 netRa11 netL11 -1.6755778754201092e-14
Rbbr11 netL11 0 80.98406978976219
Cbr11 netL11 0 -2.655614442344388e-18

* Branch 12
Rabr12 node_3 netRa12 -2.472543784195814
Lbr12 netRa12 netL12 3.518393624262684e-16
Rbbr12 netL12 0 2.5234465721550348
Cbr12 netL12 0 5.607302941093022e-17

* Branch 13
Rabr13 node_3 netRa13 1.6666091454837153
Lbr13 netRa13 netL13 3.267850105055969e-16
Rbbr13 netL13 0 -1.7329375716328606
Cbr13 netL13 0 1.1399049849777032e-16

* Branch 14
Rabr14 node_3 netRa14 -0.0013713494892064848
Lbr14 netRa14 netL14 -7.277238521870127e-17
Rbbr14 netL14 0 -4.593100533587393
Cbr14 netL14 0 -1.3416788695622425e-14

* Branch 15
Rabr15 node_3 netRa15 -0.005924348741015939
Lbr15 netRa15 netL15 1.3213111188983466e-16
Rbbr15 netL15 0 1.8584470645186466
Cbr15 netL15 0 7.353833549376253e-15

* Branch 16
Rabr16 node_3 netRa16 -716.8822125364408
Lbr16 netRa16 netL16 -3.0275617809515776e-13
Rbbr16 netL16 0 786.9792100102601
Cbr16 netL16 0 -5.424182864141664e-19

* Branch 17
Rabr17 node_3 netRa17 -199170.9921785865
Lbr17 netRa17 netL17 6.468480901258921e-12
Rbbr17 netL17 0 199298.92033916982
Cbr17 netL17 0 1.6282340089520665e-22

* Branch 18
Rabr18 node_3 netRa18 -117.24304905472633
Lbr18 netRa18 netL18 -1.2939883300550825e-13
Rbbr18 netL18 0 212.1949987735184
Cbr18 netL18 0 -5.340939445464877e-18

* Branch 19
Rabr19 node_3 netRa19 0.4226443896378112
Lbr19 netRa19 netL19 1.4040803913637558e-15
Rbbr19 netL19 0 -5.525863459282546
Cbr19 netL19 0 6.516637617119439e-16

* Branch 20
Rabr20 node_3 netRa20 -146.68633945979627
Lbr20 netRa20 netL20 8.838859520133021e-14
Rbbr20 netL20 0 202.58156685261847
Cbr20 netL20 0 2.934179184801731e-18

* Branch 21
Rabr21 node_3 netRa21 1052.2272082642944
Lbr21 netRa21 netL21 1.1144195912764549e-12
Rbbr21 netL21 0 -4064.420793698342
Cbr21 netL21 0 2.667691650513198e-19

* Branch 22
Rabr22 node_3 netRa22 1165.0928410779659
Lbr22 netRa22 netL22 -5.885575699630531e-12
Rbbr22 netL22 0 -88363.58301034331
Cbr22 netL22 0 -5.157704162140648e-20

* Branch 23
Rabr23 node_3 netRa23 1486.9379112024155
Lbr23 netRa23 netL23 1.4185714913576946e-12
Rbbr23 netL23 0 -4821.105961124356
Cbr23 netL23 0 2.01746839128014e-19

* Branch 24
Rabr24 node_3 netRa24 -14.498833775517856
Lbr24 netRa24 netL24 -3.379053855618987e-15
Rbbr24 netL24 0 16.84160357045367
Cbr24 netL24 0 -1.3898618328352756e-17

* Branch 25
Rabr25 node_3 netRa25 -93.09874542674544
Lbr25 netRa25 netL25 -2.3610096481078687e-14
Rbbr25 netL25 0 111.01240782199397
Cbr25 netL25 0 -2.2952291239958307e-18

* Branch 26
Rabr26 node_3 netRa26 2372.7804876550636
Lbr26 netRa26 netL26 1.3161804330283997e-12
Rbbr26 netL26 0 -4082.252792511775
Cbr26 netL26 0 1.3722401333849695e-19

* Branch 27
Rabr27 node_3 netRa27 -1.1385429094904063
Lbr27 netRa27 netL27 1.624078741610097e-15
Rbbr27 netL27 0 7.833078979883458
Cbr27 netL27 0 1.778270127334092e-16

* Branch 28
Rabr28 node_3 netRa28 -414.80925347854696
Lbr28 netRa28 netL28 1.3822740163624226e-13
Rbbr28 netL28 0 460.4401813248269
Cbr28 netL28 0 7.200876964755714e-19

* Branch 29
Rabr29 node_3 netRa29 150.47144522201725
Lbr29 netRa29 netL29 3.958017720569663e-14
Rbbr29 netL29 0 -161.3194715229671
Cbr29 netL29 0 1.6370078702674767e-18

* Branch 30
Rabr30 node_3 netRa30 1253.9944394020288
Lbr30 netRa30 netL30 5.257401245179587e-13
Rbbr30 netL30 0 -1882.1916212895492
Cbr30 netL30 0 2.2413927314523797e-19

* Branch 31
Rabr31 node_3 netRa31 -1115.1150749076512
Lbr31 netRa31 netL31 1.8131409994764527e-12
Rbbr31 netL31 0 8617.40049368156
Cbr31 netL31 0 1.8439888524862148e-19

* Branch 32
Rabr32 node_3 netRa32 15136.60222688622
Lbr32 netRa32 netL32 1.4412390787191742e-11
Rbbr32 netL32 0 -25138.739066589562
Cbr32 netL32 0 3.8391452768627934e-20

* Branch 33
Rabr33 node_3 netRa33 -1243.3973889089536
Lbr33 netRa33 netL33 -4.0070867151172226e-13
Rbbr33 netL33 0 1597.7298124338229
Cbr33 netL33 0 -2.025900114205754e-19

* Branch 34
Rabr34 node_3 netRa34 842.168064452698
Lbr34 netRa34 netL34 1.917334229312147e-12
Rbbr34 netL34 0 -11535.179887342667
Cbr34 netL34 0 2.036477495372627e-19

* Branch 35
Rabr35 node_3 netRa35 -515.8760415058945
Lbr35 netRa35 netL35 5.548379807247225e-13
Rbbr35 netL35 0 1780.0547425057403
Cbr35 netL35 0 5.956083654901486e-19

* Branch 36
Rabr36 node_3 netRa36 110.58944926159597
Lbr36 netRa36 netL36 6.936256500074504e-13
Rbbr36 netL36 0 -2563.0600358782112
Cbr36 netL36 0 2.6710841696637736e-18

* Branch 37
Rabr37 node_3 netRa37 -14521.319451883744
Lbr37 netRa37 netL37 1.5245033278409973e-11
Rbbr37 netL37 0 67853.28528870524
Cbr37 netL37 0 1.528221538087289e-20

* Branch 38
Rabr38 node_3 netRa38 -1570.1511544268078
Lbr38 netRa38 netL38 2.354273640842946e-12
Rbbr38 netL38 0 12341.778402977861
Cbr38 netL38 0 1.1946533432761382e-19

* Branch 39
Rabr39 node_3 netRa39 1381.942635369381
Lbr39 netRa39 netL39 9.446384072417294e-12
Rbbr39 netL39 0 -244224.20124932402
Cbr39 netL39 0 3.000260538894265e-20

* Branch 40
Rabr40 node_3 netRa40 404817.36012507597
Lbr40 netRa40 netL40 -1.0862665101386171e-10
Rbbr40 netL40 0 -428732.07828953315
Cbr40 netL40 0 -6.245441263104225e-22

* Branch 41
Rabr41 node_3 netRa41 -1437.2352193962317
Lbr41 netRa41 netL41 4.0253809229946966e-12
Rbbr41 netL41 0 30653.81252902542
Cbr41 netL41 0 8.938855874869846e-20

* Branch 42
Rabr42 node_3 netRa42 137177.2831501294
Lbr42 netRa42 netL42 8.840553063641752e-12
Rbbr42 netL42 0 -138470.9296085178
Cbr42 netL42 0 4.656473728024468e-22

* Branch 43
Rabr43 node_3 netRa43 -1515503.733588471
Lbr43 netRa43 netL43 2.394566141702164e-11
Rbbr43 netL43 0 1516664.6323591745
Cbr43 netL43 0 1.0416636532689757e-23

* Branch 44
Rabr44 node_3 netRa44 3748.020992119193
Lbr44 netRa44 netL44 1.7150308362654124e-11
Rbbr44 netL44 0 -102546.0500747401
Cbr44 netL44 0 4.611279330505103e-20

* Branch 45
Rabr45 node_3 netRa45 4038.40526656078
Lbr45 netRa45 netL45 -8.437677642139979e-12
Rbbr45 netL45 0 -23481.86878886082
Cbr45 netL45 0 -8.770456754836718e-20

* Branch 46
Rabr46 node_3 netRa46 1528.1415550537627
Lbr46 netRa46 netL46 2.2066990551483685e-13
Rbbr46 netL46 0 -1622.3000518865192
Cbr46 netL46 0 8.909606882514736e-20

* Branch 47
Rabr47 node_3 netRa47 -15.008656958216568
Lbr47 netRa47 netL47 -1.9524871683645934e-14
Rbbr47 netL47 0 85.51118202217094
Cbr47 netL47 0 -1.5339423607544788e-17

* Branch 48
Rabr48 node_3 netRa48 167.93644144537447
Lbr48 netRa48 netL48 8.579800479910934e-13
Rbbr48 netL48 0 -9639.2274171192
Cbr48 netL48 0 5.469733350627565e-19

* Branch 49
Rabr49 node_3 netRa49 5819968.837522759
Lbr49 netRa49 netL49 1.2447510144262698e-10
Rbbr49 netL49 0 -5823745.343245815
Cbr49 netL49 0 3.672953572516019e-24

* Branch 50
Rabr50 node_3 netRa50 3631.0956452431356
Lbr50 netRa50 netL50 6.995630942517391e-13
Rbbr50 netL50 0 -3849.5038540898845
Cbr50 netL50 0 5.0099544560272576e-20

* Branch 51
Rabr51 node_3 netRa51 646.5759794154104
Lbr51 netRa51 netL51 2.485038759339585e-13
Rbbr51 netL51 0 -834.456329097968
Cbr51 netL51 0 4.615224688330526e-19

* Branch 52
Rabr52 node_3 netRa52 405.1844616707883
Lbr52 netRa52 netL52 4.5085367208683456e-13
Rbbr52 netL52 0 -1419.1603341366706
Cbr52 netL52 0 7.885039452516351e-19

* Branch 53
Rabr53 node_3 netRa53 797152.8742456007
Lbr53 netRa53 netL53 -7.682560853355554e-11
Rbbr53 netL53 0 -807367.4608744315
Cbr53 netL53 0 -1.1931291102339299e-22

* Branch 54
Rabr54 node_3 netRa54 -19863.720548794994
Lbr54 netRa54 netL54 1.3143566909650295e-11
Rbbr54 netL54 0 42108.63915654514
Cbr54 netL54 0 1.566382540254579e-20

* Branch 55
Rabr55 node_3 netRa55 -376936.9089513246
Lbr55 netRa55 netL55 -1.0912206552782479e-10
Rbbr55 netL55 0 416927.5963872152
Cbr55 netL55 0 -6.952651515335154e-22

* Branch 56
Rabr56 node_3 netRa56 4567.084465368694
Lbr56 netRa56 netL56 9.392220951189875e-13
Rbbr56 netL56 0 -4998.454277246951
Cbr56 netL56 0 4.118042387347625e-20

* Branch 57
Rabr57 node_3 netRa57 356999.1768214147
Lbr57 netRa57 netL57 -7.772557758386582e-11
Rbbr57 netL57 0 -411238.67720683623
Cbr57 netL57 0 -5.289131880945706e-22

* Branch 58
Rabr58 node_3 netRa58 -372847.8180115313
Lbr58 netRa58 netL58 -9.985121944635761e-11
Rbbr58 netL58 0 407625.74993396
Cbr58 netL58 0 -6.577268271906675e-22

* Branch 59
Rabr59 node_3 netRa59 121070.0799504108
Lbr59 netRa59 netL59 9.995208952513873e-11
Rbbr59 netL59 0 -184218.98449872108
Cbr59 netL59 0 4.496207343954499e-21

* Branch 60
Rabr60 node_3 netRa60 272.4929288706348
Lbr60 netRa60 netL60 6.644635612751954e-13
Rbbr60 netL60 0 -3630.152807877534
Cbr60 netL60 0 6.781134361357738e-19

* Branch 61
Rabr61 node_3 netRa61 -339.0321550257848
Lbr61 netRa61 netL61 -4.0588328122133853e-13
Rbbr61 netL61 0 1199.3355170310579
Cbr61 netL61 0 -1.0028427350015834e-18

* Branch 62
Rabr62 node_3 netRa62 4349.530678761568
Lbr62 netRa62 netL62 -3.3041470688417156e-12
Rbbr62 netL62 0 -8275.966162898227
Cbr62 netL62 0 -9.156483059982366e-20

* Branch 63
Rabr63 node_3 netRa63 141072.41267569485
Lbr63 netRa63 netL63 9.218971691931106e-12
Rbbr63 netL63 0 -141964.01628262008
Cbr63 netL63 0 4.6041129488328495e-22

* Branch 64
Rabr64 node_3 netRa64 29229.36839720095
Lbr64 netRa64 netL64 4.278941715648979e-11
Rbbr64 netL64 0 -102203.1661977638
Cbr64 netL64 0 1.4384874318526278e-20

* Branch 65
Rabr65 node_3 netRa65 -142818.59966636205
Lbr65 netRa65 netL65 3.246146822682709e-11
Rbbr65 netL65 0 161090.46667532812
Cbr65 netL65 0 1.4100373585683585e-21

* Branch 66
Rabr66 node_3 netRa66 197280.6094789943
Lbr66 netRa66 netL66 -7.440605444422197e-11
Rbbr66 netL66 0 -234985.551413475
Cbr66 netL66 0 -1.6033643910012118e-21

* Branch 67
Rabr67 node_3 netRa67 18326.42093398585
Lbr67 netRa67 netL67 3.24286124722988e-11
Rbbr67 netL67 0 -86870.19311694361
Cbr67 netL67 0 2.0462730575302466e-20

* Branch 68
Rabr68 node_3 netRa68 -1016.408446426722
Lbr68 netRa68 netL68 -2.544791053489015e-13
Rbbr68 netL68 0 1123.2701166307795
Cbr68 netL68 0 -2.2297849171443766e-19

* Branch 69
Rabr69 node_3 netRa69 -403.5711999038736
Lbr69 netRa69 netL69 -1.6139578816325394e-13
Rbbr69 netL69 0 525.5716954793942
Cbr69 netL69 0 -7.613487856858704e-19

* Branch 70
Rabr70 node_3 netRa70 22842.62431512669
Lbr70 netRa70 netL70 5.662965243854351e-12
Rbbr70 netL70 0 -24880.08984843355
Cbr70 netL70 0 9.966664817154483e-21

* Branch 71
Rabr71 node_3 netRa71 -269.8964823042878
Lbr71 netRa71 netL71 -2.9940027803072067e-13
Rbbr71 netL71 0 867.6950426969598
Cbr71 netL71 0 -1.2795303893291996e-18

* Branch 72
Rabr72 node_3 netRa72 -10702.454623250964
Lbr72 netRa72 netL72 -1.0558316363263968e-11
Rbbr72 netL72 0 26337.665237975605
Cbr72 netL72 0 -3.7468887801142674e-20

* Branch 73
Rabr73 node_3 netRa73 16859.370404945832
Lbr73 netRa73 netL73 -5.7908211284591255e-12
Rbbr73 netL73 0 -20113.816796772324
Cbr73 netL73 0 -1.707495719509742e-20

* Branch 74
Rabr74 node_3 netRa74 -5349.961834680472
Lbr74 netRa74 netL74 -2.815580448633583e-12
Rbbr74 netL74 0 7615.412612777594
Cbr74 netL74 0 -6.910899210700288e-20

* Branch 75
Rabr75 node_3 netRa75 -4796.715133559482
Lbr75 netRa75 netL75 -2.3648789561686975e-12
Rbbr75 netL75 0 8359.962668040862
Cbr75 netL75 0 -5.897763963091063e-20

* Branch 76
Rabr76 node_3 netRa76 -4275.54493540667
Lbr76 netRa76 netL76 -2.1454024934901693e-12
Rbbr76 netL76 0 6114.173484940441
Cbr76 netL76 0 -8.208092067394105e-20

* Branch 77
Rabr77 node_3 netRa77 -150.10629308798931
Lbr77 netRa77 netL77 1.9318982295646934e-13
Rbbr77 netL77 0 702.1120311754211
Cbr77 netL77 0 1.832275234403003e-18

* Branch 78
Rabr78 node_3 netRa78 108547.11360979483
Lbr78 netRa78 netL78 -3.072930882454653e-11
Rbbr78 netL78 0 -112835.04488912484
Cbr78 netL78 0 -2.508565640445819e-21

* Branch 79
Rabr79 node_3 netRa79 -171748.93951187882
Lbr79 netRa79 netL79 4.487861605320016e-10
Rbbr79 netL79 0 1178524.248544057
Cbr79 netL79 0 2.2137041224133566e-21

* Branch 80
Rabr80 node_3 netRa80 -2229.635147469127
Lbr80 netRa80 netL80 3.2670813425429803e-12
Rbbr80 netL80 0 12712.684272047622
Cbr80 netL80 0 1.1513054391688168e-19

* Branch 81
Rabr81 node_3 netRa81 -1483849.259028696
Lbr81 netRa81 netL81 -2.339864748180237e-10
Rbbr81 netL81 0 1605699.3556154298
Cbr81 netL81 0 -9.821948575599888e-23

* Branch 82
Rabr82 node_3 netRa82 1.1628466899085101
Lbr82 netRa82 netL82 4.979865992757042e-14
Rbbr82 netL82 0 -4328.750954826106
Cbr82 netL82 0 1.0320057872154867e-17

* Branch 83
Rabr83 node_3 netRa83 -1735.0093606814778
Lbr83 netRa83 netL83 1.683370877082661e-12
Rbbr83 netL83 0 6343.528106278443
Cbr83 netL83 0 1.5279740897188155e-19

* Branch 84
Rabr84 node_3 netRa84 -16327.297513226124
Lbr84 netRa84 netL84 3.0710516947724077e-11
Rbbr84 netL84 0 57369.1317546283
Cbr84 netL84 0 3.2699280202673234e-20

* Branch 85
Rabr85 node_3 netRa85 11.266206685266352
Lbr85 netRa85 netL85 4.7633281701646795e-14
Rbbr85 netL85 0 -399.4955844591963
Cbr85 netL85 0 1.0660815611766362e-17

* Branch 86
Rabr86 node_3 netRa86 -70.02977545018422
Lbr86 netRa86 netL86 -1.4212400506698316e-13
Rbbr86 netL86 0 602.5262967695126
Cbr86 netL86 0 -3.383878502186747e-18

* Branch 87
Rabr87 node_3 netRa87 -35.082345051835674
Lbr87 netRa87 netL87 -1.0084220539248574e-13
Rbbr87 netL87 0 521.6376927492943
Cbr87 netL87 0 -5.547518176772243e-18

* Branch 88
Rabr88 node_3 netRa88 -24.38062618245233
Lbr88 netRa88 netL88 -3.7914016804517663e-14
Rbbr88 netL88 0 135.28104191902585
Cbr88 netL88 0 -1.1545053809158876e-17

* Branch 89
Rabr89 node_3 netRa89 7085.864418141988
Lbr89 netRa89 netL89 -1.936501759059948e-11
Rbbr89 netL89 0 -191096.78912408784
Cbr89 netL89 0 -1.4180252127174724e-20

* Branch 90
Rabr90 node_3 netRa90 -13925.847716650163
Lbr90 netRa90 netL90 -1.936085434646261e-11
Rbbr90 netL90 0 104644.7055928942
Cbr90 netL90 0 -1.3353950653300035e-20

* Branch 91
Rabr91 node_3 netRa91 488.48472373182386
Lbr91 netRa91 netL91 -1.5717240536538119e-12
Rbbr91 netL91 0 -2809.970423162724
Cbr91 netL91 0 -1.125423169920561e-18

* Branch 92
Rabr92 node_3 netRa92 -1419.5716771385753
Lbr92 netRa92 netL92 -1.6234920129238518e-12
Rbbr92 netL92 0 2305.2358779293495
Cbr92 netL92 0 -5.0001689802939425e-19

* Branch 93
Rabr93 node_3 netRa93 13.543300597438504
Lbr93 netRa93 netL93 1.7515459575395054e-14
Rbbr93 netL93 0 -76.4788232010023
Cbr93 netL93 0 1.70658928011929e-17

* Branch 94
Rabr94 node_3 netRa94 -7671.839556696833
Lbr94 netRa94 netL94 -2.2281121894600544e-11
Rbbr94 netL94 0 68201.98518245954
Cbr94 netL94 0 -4.4544051819213376e-20

* Branch 95
Rabr95 node_3 netRa95 23.08328549887244
Lbr95 netRa95 netL95 -3.5306754932633105e-15
Rbbr95 netL95 0 -24.67972602222607
Cbr95 netL95 0 -6.1813339752546844e-18

* Branch 96
Rabr96 node_3 netRa96 -11382.037404279285
Lbr96 netRa96 netL96 1.0628329942498157e-11
Rbbr96 netL96 0 19302.614041082816
Cbr96 netL96 0 4.7264758375106083e-20

* Branch 97
Rabr97 node_3 netRa97 19.688264457360138
Lbr97 netRa97 netL97 -2.048790859894065e-15
Rbbr97 netL97 0 -19.903817408019727
Cbr97 netL97 0 -5.202132528245554e-18

* Branch 98
Rabr98 node_3 netRa98 0.03237149667097077
Lbr98 netRa98 netL98 7.718592352964741e-17
Rbbr98 netL98 0 -0.1772760505940392
Cbr98 netL98 0 1.623126950803508e-14

* Branch 99
Rabr99 node_3 netRa99 -0.040909525712347725
Lbr99 netRa99 netL99 1.7961930129061788e-16
Rbbr99 netL99 0 0.37914602177995393
Cbr99 netL99 0 8.57007967201277e-15

.ends


* Y'34
.subckt yp34 node_3 node_4
* Branch 0
Rabr0 node_3 netRa0 4867.948183309086
Lbr0 netRa0 netL0 -2.3066826941682554e-13
Rbbr0 netL0 node_4 -4875.853370160529
Cbr0 netL0 node_4 -9.66843552833041e-21

* Branch 1
Rabr1 node_3 netRa1 2799.7476016481614
Lbr1 netRa1 netL1 -1.926205413326804e-13
Rbbr1 netL1 node_4 -2809.3707479524023
Cbr1 netL1 node_4 -2.4308394441439307e-20

* Branch 2
Rabr2 node_3 netRa2 501.93765295187364
Lbr2 netRa2 netL2 7.704859002261752e-14
Rbbr2 netL2 node_4 -510.68836011060256
Cbr2 netL2 node_4 3.054556396863629e-19

* Branch 3
Rabr3 node_3 netRa3 7.223048801665948
Lbr3 netRa3 netL3 1.6953005727917533e-14
Rbbr3 netL3 node_4 -44.0096549538837
Cbr3 netL3 node_4 6.714310442767154e-17

* Branch 4
Rabr4 node_3 netRa4 24.166271413150884
Lbr4 netRa4 netL4 3.1065331999725396e-14
Rbbr4 netL4 node_4 -44.79526135410345
Cbr4 netL4 node_4 3.0838694471577763e-17

* Branch 5
Rabr5 node_3 netRa5 4.739588208979348
Lbr5 netRa5 netL5 -3.004318612162894e-14
Rbbr5 netL5 node_4 -417.3948518050435
Cbr5 netL5 node_4 -1.1328464892462361e-17

* Branch 6
Rabr6 node_3 netRa6 -17.12598452792252
Lbr6 netRa6 netL6 1.282261353611074e-13
Rbbr6 netL6 node_4 300.0648043141687
Cbr6 netL6 node_4 1.7850834714036382e-17

* Branch 7
Rabr7 node_3 netRa7 -1.9999426126693975
Lbr7 netRa7 netL7 -3.6246787316529e-15
Rbbr7 netL7 node_4 7.5049228064113
Cbr7 netL7 node_4 -2.644851320577161e-16

* Branch 8
Rabr8 node_3 netRa8 47994.372171230716
Lbr8 netRa8 netL8 -8.31018006365199e-12
Rbbr8 netL8 node_4 -52856.3389712718
Cbr8 netL8 node_4 -3.255721382137347e-21

* Branch 9
Rabr9 node_3 netRa9 3030.5064840194887
Lbr9 netRa9 netL9 -1.820282517681046e-13
Rbbr9 netL9 node_4 -3058.626930189537
Cbr9 netL9 node_4 -1.9600484934853588e-20

* Branch 10
Rabr10 node_3 netRa10 64.94586542922522
Lbr10 netRa10 netL10 -2.6960808225386837e-14
Rbbr10 netL10 node_4 -94.87752571257928
Cbr10 netL10 node_4 -4.319708567805439e-18

* Branch 11
Rabr11 node_3 netRa11 12.35260168278153
Lbr11 netRa11 netL11 2.0806733866269074e-14
Rbbr11 netL11 node_4 -94.04896631646045
Cbr11 netL11 node_4 1.879628691466752e-17

* Branch 12
Rabr12 node_3 netRa12 181.2266483827361
Lbr12 netRa12 netL12 5.694834611901528e-14
Rbbr12 netL12 node_4 -225.0653213114128
Cbr12 netL12 node_4 1.4085637264514446e-18

* Branch 13
Rabr13 node_3 netRa13 2458.1734924300704
Lbr13 netRa13 netL13 3.0617642704888115e-12
Rbbr13 netL13 node_4 -15393.387406449308
Cbr13 netL13 node_4 8.363117560645485e-20

* Branch 14
Rabr14 node_3 netRa14 352.31846328934506
Lbr14 netRa14 netL14 6.56494852538522e-14
Rbbr14 netL14 node_4 -380.1154958731277
Cbr14 netL14 node_4 4.925829232782718e-19

* Branch 15
Rabr15 node_3 netRa15 -1758.0994865263847
Lbr15 netRa15 netL15 2.0873417847882156e-13
Rbbr15 netL15 node_4 1832.6720906463102
Cbr15 netL15 node_4 6.458654021942481e-20

* Branch 16
Rabr16 node_3 netRa16 -7.7762295868836055
Lbr16 netRa16 netL16 9.424549556324194e-14
Rbbr16 netL16 node_4 2645.3597695502626
Cbr16 netL16 node_4 3.512178235164217e-18

* Branch 17
Rabr17 node_3 netRa17 10.2945474191248
Lbr17 netRa17 netL17 1.1000678219319197e-14
Rbbr17 netL17 node_4 -35.88737198182563
Cbr17 netL17 node_4 3.057614059200335e-17

* Branch 18
Rabr18 node_3 netRa18 114.47226496704864
Lbr18 netRa18 netL18 -5.609125012961563e-14
Rbbr18 netL18 node_4 -196.0962729773363
Cbr18 netL18 node_4 -2.4694806077294253e-18

* Branch 19
Rabr19 node_3 netRa19 -19.89533391130622
Lbr19 netRa19 netL19 2.7941341712921864e-14
Rbbr19 netL19 node_4 89.85826604896414
Cbr19 netL19 node_4 1.5129219902334263e-17

* Branch 20
Rabr20 node_3 netRa20 43.995605696087814
Lbr20 netRa20 netL20 6.011536235066096e-14
Rbbr20 netL20 node_4 -302.10820189700587
Cbr20 netL20 node_4 4.664342075584694e-18

* Branch 21
Rabr21 node_3 netRa21 -76.0161495174671
Lbr21 netRa21 netL21 -4.485700668692898e-14
Rbbr21 netL21 node_4 105.19306743510575
Cbr21 netL21 node_4 -5.682264789491714e-18

* Branch 22
Rabr22 node_3 netRa22 -3.297053682723883
Lbr22 netRa22 netL22 3.110735972937173e-14
Rbbr22 netL22 node_4 491.93584280254925
Cbr22 netL22 node_4 1.6024604766931134e-17

* Branch 23
Rabr23 node_3 netRa23 -648.0389214148844
Lbr23 netRa23 netL23 1.121644902860195e-13
Rbbr23 netL23 node_4 676.5068521695794
Cbr23 netL23 node_4 2.5493659085456177e-19

* Branch 24
Rabr24 node_3 netRa24 -6.154937560918024
Lbr24 netRa24 netL24 3.026649695156881e-14
Rbbr24 netL24 node_4 269.8386914621649
Cbr24 netL24 node_4 1.655066667990237e-17

* Branch 25
Rabr25 node_3 netRa25 -16.569501415179914
Lbr25 netRa25 netL25 2.626076884102574e-14
Rbbr25 netL25 node_4 93.60926843532509
Cbr25 netL25 node_4 1.639757879049268e-17

* Branch 26
Rabr26 node_3 netRa26 -5.935100963929206
Lbr26 netRa26 netL26 -8.982849862142932e-14
Rbbr26 netL26 node_4 1389.7853068231498
Cbr26 netL26 node_4 -1.5739417839335687e-17

* Branch 27
Rabr27 node_3 netRa27 172.76666403052857
Lbr27 netRa27 netL27 7.17471504552196e-14
Rbbr27 netL27 node_4 -237.83356001545027
Cbr27 netL27 node_4 1.7608465655665573e-18

* Branch 28
Rabr28 node_3 netRa28 42.647924116678055
Lbr28 netRa28 netL28 4.0478450444979957e-13
Rbbr28 netL28 node_4 -14756.491104600163
Cbr28 netL28 node_4 7.931958486982389e-19

* Branch 29
Rabr29 node_3 netRa29 384.5035724074826
Lbr29 netRa29 netL29 1.47801349823035e-13
Rbbr29 netL29 node_4 -520.4815231703749
Cbr29 netL29 node_4 7.442093620679484e-19

* Branch 30
Rabr30 node_3 netRa30 8787.003753977951
Lbr30 netRa30 netL30 5.872099925095922e-13
Rbbr30 netL30 node_4 -8878.407586552514
Cbr30 netL30 node_4 7.536797961723659e-21

* Branch 31
Rabr31 node_3 netRa31 -5749.857427737778
Lbr31 netRa31 netL31 -3.4587977041417017e-13
Rbbr31 netL31 node_4 5779.770214840992
Cbr31 netL31 node_4 -1.0419780071543241e-20

* Branch 32
Rabr32 node_3 netRa32 -11.63190838354257
Lbr32 netRa32 netL32 -3.443355107558009e-14
Rbbr32 netL32 node_4 126.45511234120158
Cbr32 netL32 node_4 -2.4805054166076906e-17

* Branch 33
Rabr33 node_3 netRa33 -25.683303668038057
Lbr33 netRa33 netL33 -4.433862381731428e-14
Rbbr33 netL33 node_4 107.10707895236146
Cbr33 netL33 node_4 -1.6637127557221573e-17

* Branch 34
Rabr34 node_3 netRa34 157.57089682072188
Lbr34 netRa34 netL34 -1.0122079755542059e-13
Rbbr34 netL34 node_4 -204.9082370977954
Cbr34 netL34 node_4 -3.099267790722226e-18

* Branch 35
Rabr35 node_3 netRa35 98.24129339466785
Lbr35 netRa35 netL35 -1.1163458960526623e-13
Rbbr35 netL35 node_4 -423.9756361773948
Cbr35 netL35 node_4 -2.626952914284883e-18

* Branch 36
Rabr36 node_3 netRa36 -537.5765901821799
Lbr36 netRa36 netL36 -1.4392949519656141e-13
Rbbr36 netL36 node_4 580.888852637013
Cbr36 netL36 node_4 -4.630998214908643e-19

* Branch 37
Rabr37 node_3 netRa37 -29854.893463748434
Lbr37 netRa37 netL37 1.0037029489238444e-12
Rbbr37 netL37 node_4 29882.429974895786
Cbr37 netL37 node_4 1.1244060159989354e-21

* Branch 38
Rabr38 node_3 netRa38 -131.28615101234448
Lbr38 netRa38 netL38 -9.601310053913055e-14
Rbbr38 netL38 node_4 195.07392398838405
Cbr38 netL38 node_4 -3.794587981284372e-18

* Branch 39
Rabr39 node_3 netRa39 -13.28738622515219
Lbr39 netRa39 netL39 2.4427807734278386e-14
Rbbr39 netL39 node_4 88.63451006723514
Cbr39 netL39 node_4 2.0149608186542273e-17

* Branch 40
Rabr40 node_3 netRa40 -1716.847181661214
Lbr40 netRa40 netL40 2.094674078882516e-13
Rbbr40 netL40 node_4 1756.911547606928
Cbr40 netL40 node_4 6.930962179621091e-20

* Branch 41
Rabr41 node_3 netRa41 -18.81563297065073
Lbr41 netRa41 netL41 3.8029121928558273e-14
Rbbr41 netL41 node_4 150.3026660498265
Cbr41 netL41 node_4 1.3033984926349041e-17

* Branch 42
Rabr42 node_3 netRa42 -75.95091286889998
Lbr42 netRa42 netL42 -8.63062193469827e-14
Rbbr42 netL42 node_4 168.5151428828518
Cbr42 netL42 node_4 -6.863513508634183e-18

* Branch 43
Rabr43 node_3 netRa43 -2320.4206790290123
Lbr43 netRa43 netL43 -2.4084217389749295e-13
Rbbr43 netL43 node_4 2355.483115401712
Cbr43 netL43 node_4 -4.41337432575429e-20

* Branch 44
Rabr44 node_3 netRa44 48.492940106853176
Lbr44 netRa44 netL44 -1.1180354829097865e-13
Rbbr44 netL44 node_4 -658.4892508920439
Cbr44 netL44 node_4 -3.383069125575192e-18

* Branch 45
Rabr45 node_3 netRa45 -38.59349290611335
Lbr45 netRa45 netL45 5.5725313167880346e-14
Rbbr45 netL45 node_4 180.47787398571725
Cbr45 netL45 node_4 7.82911588635638e-18

* Branch 46
Rabr46 node_3 netRa46 -1390.4763832910526
Lbr46 netRa46 netL46 -1.4942939551482728e-13
Rbbr46 netL46 node_4 1416.4114870196006
Cbr46 netL46 node_4 -7.599560007551984e-20

* Branch 47
Rabr47 node_3 netRa47 -1557.1085121121944
Lbr47 netRa47 netL47 -2.940590551071088e-13
Rbbr47 netL47 node_4 1604.1070991837923
Cbr47 netL47 node_4 -1.1806247416676396e-19

* Branch 48
Rabr48 node_3 netRa48 58.70398515703119
Lbr48 netRa48 netL48 4.8664097869583336e-14
Rbbr48 netL48 node_4 -162.35730342565944
Cbr48 netL48 node_4 5.168412687241137e-18

* Branch 49
Rabr49 node_3 netRa49 -194.04435610636642
Lbr49 netRa49 netL49 -1.2951026925216838e-13
Rbbr49 netL49 node_4 270.0469295915964
Cbr49 netL49 node_4 -2.4936421615904653e-18

* Branch 50
Rabr50 node_3 netRa50 -5350.361890800546
Lbr50 netRa50 netL50 -3.8403546752100783e-13
Rbbr50 netL50 node_4 5392.040466707516
Cbr50 netL50 node_4 -1.3324423521975482e-20

* Branch 51
Rabr51 node_3 netRa51 -34.36640287412781
Lbr51 netRa51 netL51 -5.2808413226759575e-14
Rbbr51 netL51 node_4 117.20396324629483
Cbr51 netL51 node_4 -1.3372671861000617e-17

* Branch 52
Rabr52 node_3 netRa52 -141.99857485908692
Lbr52 netRa52 netL52 5.2546164478841735e-14
Rbbr52 netL52 node_4 182.69716453829545
Cbr52 netL52 node_4 2.015969699921842e-18

* Branch 53
Rabr53 node_3 netRa53 -65.286584733514
Lbr53 netRa53 netL53 7.473158292574778e-14
Rbbr53 netL53 node_4 237.12600206119893
Cbr53 netL53 node_4 4.76223743418296e-18

* Branch 54
Rabr54 node_3 netRa54 -31.947324750668656
Lbr54 netRa54 netL54 -8.290195394712423e-14
Rbbr54 netL54 node_4 244.06617671989483
Cbr54 netL54 node_4 -1.0953928985559338e-17

* Branch 55
Rabr55 node_3 netRa55 -78.78825498531069
Lbr55 netRa55 netL55 5.0097803737934204e-14
Rbbr55 netL55 node_4 132.51599055012616
Cbr55 netL55 node_4 4.76544672933137e-18

* Branch 56
Rabr56 node_3 netRa56 -177.0517677988171
Lbr56 netRa56 netL56 -1.1944915091138325e-13
Rbbr56 netL56 node_4 270.5484977363973
Cbr56 netL56 node_4 -2.5114860531214623e-18

* Branch 57
Rabr57 node_3 netRa57 -664.4609504497339
Lbr57 netRa57 netL57 2.380658399223725e-13
Rbbr57 netL57 node_4 824.6064699839135
Cbr57 netL57 node_4 4.3295354603531775e-19

* Branch 58
Rabr58 node_3 netRa58 -491.432704510921
Lbr58 netRa58 netL58 2.193364958794815e-13
Rbbr58 netL58 node_4 754.3327268712704
Cbr58 netL58 node_4 5.890929095036769e-19

* Branch 59
Rabr59 node_3 netRa59 -253.70895416985744
Lbr59 netRa59 netL59 1.3863073660173874e-13
Rbbr59 netL59 node_4 313.3211001083301
Cbr59 netL59 node_4 1.734737738334616e-18

* Branch 60
Rabr60 node_3 netRa60 -22724.79035294957
Lbr60 netRa60 netL60 -1.3534053896329613e-12
Rbbr60 netL60 node_4 22945.50309218445
Cbr60 netL60 node_4 -2.5969871117541555e-21

* Branch 61
Rabr61 node_3 netRa61 -75.6351745266586
Lbr61 netRa61 netL61 5.2471816280547076e-14
Rbbr61 netL61 node_4 134.83521964981873
Cbr61 netL61 node_4 5.113336917665279e-18

* Branch 62
Rabr62 node_3 netRa62 -132.93670756774432
Lbr62 netRa62 netL62 9.603696293139754e-14
Rbbr62 netL62 node_4 238.6654934180559
Cbr62 netL62 node_4 3.0080130541104496e-18

* Branch 63
Rabr63 node_3 netRa63 -20891.8290558178
Lbr63 netRa63 netL63 1.2647037886271893e-12
Rbbr63 netL63 node_4 21085.10758061141
Cbr63 netL63 node_4 2.869540064125846e-21

* Branch 64
Rabr64 node_3 netRa64 -64.87166378190945
Lbr64 netRa64 netL64 -5.3266818843939264e-14
Rbbr64 netL64 node_4 119.29397659940261
Cbr64 netL64 node_4 -6.9298404583210565e-18

* Branch 65
Rabr65 node_3 netRa65 -11026.467284847236
Lbr65 netRa65 netL65 -6.758206918038767e-13
Rbbr65 netL65 node_4 11083.20460671236
Cbr65 netL65 node_4 -5.532809991467992e-21

* Branch 66
Rabr66 node_3 netRa66 -220.04903330034614
Lbr66 netRa66 netL66 1.171489974543637e-13
Rbbr66 netL66 node_4 348.71930438474686
Cbr66 netL66 node_4 1.520192077623559e-18

* Branch 67
Rabr67 node_3 netRa67 -54.692630622459816
Lbr67 netRa67 netL67 5.410779345722595e-14
Rbbr67 netL67 node_4 143.16839800366526
Cbr67 netL67 node_4 6.856318832969025e-18

* Branch 68
Rabr68 node_3 netRa68 -7.905158749484168
Lbr68 netRa68 netL68 1.0104324277829147e-13
Rbbr68 netL68 node_4 909.4557845357698
Cbr68 netL68 node_4 1.2800974408517888e-17

* Branch 69
Rabr69 node_3 netRa69 284.9788038985007
Lbr69 netRa69 netL69 -2.5787322849340666e-13
Rbbr69 netL69 node_4 -813.9446731433186
Cbr69 netL69 node_4 -1.1040981378090763e-18

* Branch 70
Rabr70 node_3 netRa70 73.66760766722719
Lbr70 netRa70 netL70 -2.8786830942654495e-13
Rbbr70 netL70 node_4 -3122.1914653057
Cbr70 netL70 node_4 -1.2153897049981134e-18

* Branch 71
Rabr71 node_3 netRa71 -69.80615835843005
Lbr71 netRa71 netL71 -6.252536888510731e-14
Rbbr71 netL71 node_4 137.87500651738247
Cbr71 netL71 node_4 -6.540510711372479e-18

* Branch 72
Rabr72 node_3 netRa72 -12034.271789462942
Lbr72 netRa72 netL72 -3.3667517826335516e-12
Rbbr72 netL72 node_4 15264.407009941888
Cbr72 netL72 node_4 -1.8365686089109793e-20

* Branch 73
Rabr73 node_3 netRa73 2.4245961484512533
Lbr73 netRa73 netL73 -7.924828985913251e-14
Rbbr73 netL73 node_4 -2069.8479078101695
Cbr73 netL73 node_4 -1.2821421770766415e-17

* Branch 74
Rabr74 node_3 netRa74 -86.34574628929454
Lbr74 netRa74 netL74 -9.025145567454867e-14
Rbbr74 netL74 node_4 198.59958271222413
Cbr74 netL74 node_4 -5.301486282784914e-18

* Branch 75
Rabr75 node_3 netRa75 -6012.558569111008
Lbr75 netRa75 netL75 3.3194448130592013e-12
Rbbr75 netL75 node_4 11788.99542572283
Cbr75 netL75 node_4 4.665614388499882e-20

* Branch 76
Rabr76 node_3 netRa76 740.2607112306767
Lbr76 netRa76 netL76 -9.714030288089056e-13
Rbbr76 netL76 node_4 -4364.915257124543
Cbr76 netL76 node_4 -2.980624915158673e-19

* Branch 77
Rabr77 node_3 netRa77 2749.854471215716
Lbr77 netRa77 netL77 2.3791906059886455e-12
Rbbr77 netL77 node_4 -9436.664112145236
Cbr77 netL77 node_4 9.218127995955325e-20

* Branch 78
Rabr78 node_3 netRa78 -32.16918208004931
Lbr78 netRa78 netL78 -3.7204731577085776e-14
Rbbr78 netL78 node_4 87.13101015087803
Cbr78 netL78 node_4 -1.3367486616075589e-17

* Branch 79
Rabr79 node_3 netRa79 -20567.863134280044
Lbr79 netRa79 netL79 4.449277077246134e-12
Rbbr79 netL79 node_4 21210.30677620322
Cbr79 netL79 node_4 1.0187154501387615e-20

* Branch 80
Rabr80 node_3 netRa80 8987.416648729188
Lbr80 netRa80 netL80 3.4544210165225437e-12
Rbbr80 netL80 node_4 -9771.906567925447
Cbr80 netL80 node_4 3.9409917104355247e-20

* Branch 81
Rabr81 node_3 netRa81 -240.60831352913482
Lbr81 netRa81 netL81 -6.459712984156021e-13
Rbbr81 netL81 node_4 5206.57325472921
Cbr81 netL81 node_4 -5.221746055699219e-19

* Branch 82
Rabr82 node_3 netRa82 -45084.18142546388
Lbr82 netRa82 netL82 3.8066374246228785e-12
Rbbr82 netL82 node_4 46251.76974882663
Cbr82 netL82 node_4 1.8249375762194013e-21

* Branch 83
Rabr83 node_3 netRa83 -33.48092407153672
Lbr83 netRa83 netL83 -2.9163920521979126e-14
Rbbr83 netL83 node_4 66.43542824119666
Cbr83 netL83 node_4 -1.3152578830157403e-17

* Branch 84
Rabr84 node_3 netRa84 -533.3775870452743
Lbr84 netRa84 netL84 1.0588608225517226e-12
Rbbr84 netL84 node_4 1871.0031104307816
Cbr84 netL84 node_4 1.054094216360939e-18

* Branch 85
Rabr85 node_3 netRa85 1083.9793255498566
Lbr85 netRa85 netL85 2.1698947805480656e-12
Rbbr85 netL85 node_4 -3757.582278820703
Cbr85 netL85 node_4 5.358707727297785e-19

* Branch 86
Rabr86 node_3 netRa86 -187.87925010431113
Lbr86 netRa86 netL86 1.22228376280552e-13
Rbbr86 netL86 node_4 294.0981926935731
Cbr86 netL86 node_4 2.2080675050094427e-18

* Branch 87
Rabr87 node_3 netRa87 45506.683212537275
Lbr87 netRa87 netL87 -1.011871555556845e-11
Rbbr87 netL87 node_4 -46785.08543361244
Cbr87 netL87 node_4 -4.750102779721219e-21

* Branch 88
Rabr88 node_3 netRa88 3263.0146845474546
Lbr88 netRa88 netL88 2.9872999453883715e-12
Rbbr88 netL88 node_4 -12034.039788847016
Cbr88 netL88 node_4 7.624537918441666e-20

* Branch 89
Rabr89 node_3 netRa89 135.3725410441513
Lbr89 netRa89 netL89 -7.756725839948254e-13
Rbbr89 netL89 node_4 -2370.8961611516474
Cbr89 netL89 node_4 -2.385497070976926e-18

* Branch 90
Rabr90 node_3 netRa90 -35.81507512731694
Lbr90 netRa90 netL90 -6.176104117829342e-13
Rbbr90 netL90 node_4 5478.910127390079
Cbr90 netL90 node_4 -3.2763782580136928e-18

* Branch 91
Rabr91 node_3 netRa91 -51.99890201363572
Lbr91 netRa91 netL91 -5.044022359981901e-14
Rbbr91 netL91 node_4 116.46011849660887
Cbr91 netL91 node_4 -8.344294899080082e-18

* Branch 92
Rabr92 node_3 netRa92 352.9429961143817
Lbr92 netRa92 netL92 -1.6206759713701758e-12
Rbbr92 netL92 node_4 -4262.277275768444
Cbr92 netL92 node_4 -1.0708359975049667e-18

* Branch 93
Rabr93 node_3 netRa93 -293.05117028518174
Lbr93 netRa93 netL93 -7.196204602776654e-13
Rbbr93 netL93 node_4 1129.6801452881339
Cbr93 netL93 node_4 -2.1785132043698806e-18

* Branch 94
Rabr94 node_3 netRa94 1836.2233022555165
Lbr94 netRa94 netL94 -4.710520138570051e-12
Rbbr94 netL94 node_4 -8448.83935181987
Cbr94 netL94 node_4 -3.0310066629116935e-19

* Branch 95
Rabr95 node_3 netRa95 -141.46760268470783
Lbr95 netRa95 netL95 -3.448281494686965e-13
Rbbr95 netL95 node_4 518.3546593196231
Cbr95 netL95 node_4 -4.703848835398286e-18

* Branch 96
Rabr96 node_3 netRa96 -3730.7037890402216
Lbr96 netRa96 netL96 1.1598587887179198e-12
Rbbr96 netL96 node_4 3894.6147179370705
Cbr96 netL96 node_4 7.973137834100271e-20

* Branch 97
Rabr97 node_3 netRa97 3471.249047857131
Lbr97 netRa97 netL97 2.530872596278443e-12
Rbbr97 netL97 node_4 -9836.78567601796
Cbr97 netL97 node_4 7.440136167544658e-20

* Branch 98
Rabr98 node_3 netRa98 -76.73882629277973
Lbr98 netRa98 netL98 -4.385391000561237e-14
Rbbr98 netL98 node_4 153.8818839678509
Cbr98 netL98 node_4 -3.776289184416809e-18

* Branch 99
Rabr99 node_3 netRa99 105.2238078594357
Lbr99 netRa99 netL99 -3.337157735833214e-14
Rbbr99 netL99 node_4 -112.63491522489882
Cbr99 netL99 node_4 -2.715321613409974e-18

.ends


* Y'44
.subckt yp44 node_4 0
* Branch 0
Rabr0 node_4 netRa0 1309.999677498572
Lbr0 netRa0 netL0 -9.7382270823973e-14
Rbbr0 netL0 0 -1318.86742029454
Cbr0 netL0 0 -5.576336156595904e-20

* Branch 1
Rabr1 node_4 netRa1 48.22375417442098
Lbr1 netRa1 netL1 2.8188299137966655e-14
Rbbr1 netL1 0 -70.3764189744114
Cbr1 netL1 0 9.011287030566434e-18

* Branch 2
Rabr2 node_4 netRa2 -8284.081809208003
Lbr2 netRa2 netL2 -1.7064347158079838e-12
Rbbr2 netL2 0 8736.54560944088
Cbr2 netL2 0 -2.424547264816085e-20

* Branch 3
Rabr3 node_4 netRa3 -0.1508905104822364
Lbr3 netRa3 netL3 1.5724000083729218e-14
Rbbr3 netL3 0 154.94911075906117
Cbr3 netL3 0 5.136214957690692e-17

* Branch 4
Rabr4 node_4 netRa4 -15472.513303262946
Lbr4 netRa4 netL4 -1.022544133719447e-12
Rbbr4 netL4 0 15556.545985050443
Cbr4 netL4 0 -4.275879037031589e-21

* Branch 5
Rabr5 node_4 netRa5 -0.08835303039734219
Lbr5 netRa5 netL5 -4.732427846054894e-15
Rbbr5 netL5 0 -110.33656792339758
Cbr5 netL5 0 -1.7155699438625502e-16

* Branch 6
Rabr6 node_4 netRa6 3.2144591823061375
Lbr6 netRa6 netL6 2.8502279957078064e-14
Rbbr6 netL6 0 -465.63523353880925
Cbr6 netL6 0 2.900290215644367e-17

* Branch 7
Rabr7 node_4 netRa7 1.7096136058261298
Lbr7 netRa7 netL7 2.94732006819056e-14
Rbbr7 netL7 0 -1778.8266684599134
Cbr7 netL7 0 2.7198995651768644e-17

* Branch 8
Rabr8 node_4 netRa8 -175.73997763552802
Lbr8 netRa8 netL8 4.1103976267331307e-13
Rbbr8 netL8 0 1338.2438790706617
Cbr8 netL8 0 1.6397265619236734e-18

* Branch 9
Rabr9 node_4 netRa9 43.68183201578586
Lbr9 netRa9 netL9 2.0078804776089297e-14
Rbbr9 netL9 0 -69.66804275473257
Cbr9 netL9 0 6.670365695943324e-18

* Branch 10
Rabr10 node_4 netRa10 -39.25374065146807
Lbr10 netRa10 netL10 -1.5124239952080862e-14
Rbbr10 netL10 0 55.60307855437368
Cbr10 netL10 0 -6.98616565779125e-18

* Branch 11
Rabr11 node_4 netRa11 -7505.5154345115725
Lbr11 netRa11 netL11 -1.1634897942085673e-11
Rbbr11 netL11 0 61926.23291213008
Cbr11 netL11 0 -2.5809306590728557e-20

* Branch 12
Rabr12 node_4 netRa12 -122236.61503555112
Lbr12 netRa12 netL12 5.441182271784732e-11
Rbbr12 netL12 0 185118.99645984947
Cbr12 netL12 0 2.3840318684215423e-21

* Branch 13
Rabr13 node_4 netRa13 -4657.487504718507
Lbr13 netRa13 netL13 1.6220988927924406e-12
Rbbr13 netL13 0 6453.009103599979
Cbr13 netL13 0 5.362154677396502e-20

* Branch 14
Rabr14 node_4 netRa14 -378839.96052533906
Lbr14 netRa14 netL14 5.6710551378271463e-11
Rbbr14 netL14 0 394658.00979214197
Cbr14 netL14 0 3.78245109998816e-22

* Branch 15
Rabr15 node_4 netRa15 -12577.118532844355
Lbr15 netRa15 netL15 5.692015677525228e-13
Rbbr15 netL15 0 12648.644289811426
Cbr15 netL15 0 3.575089669752458e-21

* Branch 16
Rabr16 node_4 netRa16 938.7976508824299
Lbr16 netRa16 netL16 1.3430929539413708e-12
Rbbr16 netL16 0 -3196.4260114245126
Cbr16 netL16 0 4.591955871578132e-19

* Branch 17
Rabr17 node_4 netRa17 -24024.769251931713
Lbr17 netRa17 netL17 2.37566448666064e-11
Rbbr17 netL17 0 80569.02099133078
Cbr17 netL17 0 1.2076144884541605e-20

* Branch 18
Rabr18 node_4 netRa18 -27119.66155633352
Lbr18 netRa18 netL18 6.29105499407992e-13
Rbbr18 netL18 0 27148.636584980246
Cbr18 netL18 0 8.541341745391723e-22

* Branch 19
Rabr19 node_4 netRa19 -138.57996228977848
Lbr19 netRa19 netL19 8.12441774156913e-13
Rbbr19 netL19 0 13871.49105879825
Cbr19 netL19 0 3.8694106848162147e-19

* Branch 20
Rabr20 node_4 netRa20 1369.9446681866084
Lbr20 netRa20 netL20 -7.049789072837585e-13
Rbbr20 netL20 0 -2079.4450918768466
Cbr20 netL20 0 -2.4573340547146524e-19

* Branch 21
Rabr21 node_4 netRa21 1706.5547496224924
Lbr21 netRa21 netL21 -1.976593137762894e-12
Rbbr21 netL21 0 -4895.8537932754125
Cbr21 netL21 0 -2.3289623743247813e-19

* Branch 22
Rabr22 node_4 netRa22 523.8860887955428
Lbr22 netRa22 netL22 -4.778862978342328e-13
Rbbr22 netL22 0 -1888.164434270411
Cbr22 netL22 0 -4.771809985373491e-19

* Branch 23
Rabr23 node_4 netRa23 41368.584073777274
Lbr23 netRa23 netL23 3.536590815722854e-11
Rbbr23 netL23 0 -113916.23421360634
Cbr23 netL23 0 7.590518189531035e-21

* Branch 24
Rabr24 node_4 netRa24 13.124361350647524
Lbr24 netRa24 netL24 -6.441818493929214e-14
Rbbr24 netL24 0 -601.63386309286
Cbr24 netL24 0 -7.660542973164284e-18

* Branch 25
Rabr25 node_4 netRa25 6491.447356489945
Lbr25 netRa25 netL25 1.5575564901466016e-12
Rbbr25 netL25 0 -7341.603387678654
Cbr25 netL25 0 3.278471070119042e-20

* Branch 26
Rabr26 node_4 netRa26 -19669.104260290445
Lbr26 netRa26 netL26 2.8406307710709246e-11
Rbbr26 netL26 0 89260.29539445172
Cbr26 netL26 0 1.588253080147026e-20

* Branch 27
Rabr27 node_4 netRa27 9753.262800428221
Lbr27 netRa27 netL27 -8.314161329597658e-12
Rbbr27 netL27 0 -19261.346493682795
Cbr27 netL27 0 -4.3798021928440095e-20

* Branch 28
Rabr28 node_4 netRa28 -208.2231268606269
Lbr28 netRa28 netL28 -1.8229397762929634e-13
Rbbr28 netL28 0 571.9326027580779
Cbr28 netL28 0 -1.5466876780579212e-18

* Branch 29
Rabr29 node_4 netRa29 -15730.624400185787
Lbr29 netRa29 netL29 1.5649455817752035e-12
Rbbr29 netL29 0 16160.851967094795
Cbr29 netL29 0 6.148933563643991e-21

* Branch 30
Rabr30 node_4 netRa30 16912517.254040234
Lbr30 netRa30 netL30 -2.6724970717984085e-09
Rbbr30 netL30 0 -17283694.50909342
Cbr30 netL30 0 -9.126476200311032e-24

* Branch 31
Rabr31 node_4 netRa31 2568.1305005391187
Lbr31 netRa31 netL31 2.9695557578339437e-12
Rbbr31 netL31 0 -6442.528814141438
Cbr31 netL31 0 1.8180959129410366e-19

* Branch 32
Rabr32 node_4 netRa32 1010626.9124903692
Lbr32 netRa32 netL32 1.0054976040005639e-10
Rbbr32 netL32 0 -1033822.8672349309
Cbr32 netL32 0 9.634171888963373e-23

* Branch 33
Rabr33 node_4 netRa33 -273470.6938702417
Lbr33 netRa33 netL33 1.9701466980688088e-09
Rbbr33 netL33 0 11481664.311698044
Cbr33 netL33 0 5.825125476280247e-22

* Branch 34
Rabr34 node_4 netRa34 21236.167384431712
Lbr34 netRa34 netL34 -6.37654201722072e-11
Rbbr34 netL34 0 -169308.71512004707
Cbr34 netL34 0 -1.7215925530399115e-20

* Branch 35
Rabr35 node_4 netRa35 -17992.182617169517
Lbr35 netRa35 netL35 -8.157058047306071e-11
Rbbr35 netL35 0 300425.28962241905
Cbr35 netL35 0 -1.575339500303344e-20

* Branch 36
Rabr36 node_4 netRa36 -1815.408024037834
Lbr36 netRa36 netL36 -4.362036001087737e-12
Rbbr36 netL36 0 25079.575335173264
Cbr36 netL36 0 -9.784896794545033e-20

* Branch 37
Rabr37 node_4 netRa37 500.18563470462584
Lbr37 netRa37 netL37 1.1551975114874053e-12
Rbbr37 netL37 0 -8144.308732002012
Cbr37 netL37 0 2.8905595994263005e-19

* Branch 38
Rabr38 node_4 netRa38 -17917.274138639095
Lbr38 netRa38 netL38 -4.821376114856442e-11
Rbbr38 netL38 0 108619.98476759369
Cbr38 netL38 0 -2.5331896372177663e-20

* Branch 39
Rabr39 node_4 netRa39 5643810.002350252
Lbr39 netRa39 netL39 1.3717622723076551e-10
Rbbr39 netL39 0 -5648450.638111455
Cbr39 netL39 0 4.3038985976560985e-24

* Branch 40
Rabr40 node_4 netRa40 -7296.867947660223
Lbr40 netRa40 netL40 -4.2506713585155455e-11
Rbbr40 netL40 0 264451.47888641007
Cbr40 netL40 0 -2.3088288113276317e-20

* Branch 41
Rabr41 node_4 netRa41 5380.077315948166
Lbr41 netRa41 netL41 -1.2726358961741527e-10
Rbbr41 netL41 0 -1806340.6361709016
Cbr41 netL41 0 -1.1206509429121668e-20

* Branch 42
Rabr42 node_4 netRa42 -12048261.951731637
Lbr42 netRa42 netL42 -1.2145556704514424e-09
Rbbr42 netL42 0 12149648.605767649
Cbr42 netL42 0 -8.303063919814731e-24

* Branch 43
Rabr43 node_4 netRa43 -17648.891340508242
Lbr43 netRa43 netL43 -3.211904368009046e-11
Rbbr43 netL43 0 222174.54035444956
Cbr43 netL43 0 -8.29606543219498e-21

* Branch 44
Rabr44 node_4 netRa44 9262.967449842447
Lbr44 netRa44 netL44 -3.0369049179274007e-12
Rbbr44 netL44 0 -10455.994866786437
Cbr44 netL44 0 -3.129306632556753e-20

* Branch 45
Rabr45 node_4 netRa45 -109281.09136160168
Lbr45 netRa45 netL45 -2.6246633980477732e-11
Rbbr45 netL45 0 118326.7967205685
Cbr45 netL45 0 -2.032623279336124e-21

* Branch 46
Rabr46 node_4 netRa46 -12730.713458703774
Lbr46 netRa46 netL46 -3.8286346923535084e-11
Rbbr46 netL46 0 125857.66487358666
Cbr46 netL46 0 -2.4321621469071955e-20

* Branch 47
Rabr47 node_4 netRa47 -8989.227200828975
Lbr47 netRa47 netL47 -4.0572363168750954e-11
Rbbr47 netL47 0 132994.61669379307
Cbr47 netL47 0 -3.483942138490075e-20

* Branch 48
Rabr48 node_4 netRa48 139.10300470900302
Lbr48 netRa48 netL48 -1.7128159614338873e-11
Rbbr48 netL48 0 -2628364.0277338624
Cbr48 netL48 0 -2.7479263076245795e-20

* Branch 49
Rabr49 node_4 netRa49 -4871.803776408088
Lbr49 netRa49 netL49 8.841565413002971e-12
Rbbr49 netL49 0 22314.322057155474
Cbr49 netL49 0 8.050684286752162e-20

* Branch 50
Rabr50 node_4 netRa50 6461.669980869315
Lbr50 netRa50 netL50 1.15930406320456e-11
Rbbr50 netL50 0 -41385.61602932977
Cbr50 netL50 0 4.378956490847723e-20

* Branch 51
Rabr51 node_4 netRa51 -1368814.444927805
Lbr51 netRa51 netL51 -2.5929048167459335e-10
Rbbr51 netL51 0 1494534.9431912377
Cbr51 netL51 0 -1.2687622550820772e-22

* Branch 52
Rabr52 node_4 netRa52 -102712764.07129928
Lbr52 netRa52 netL52 -1.6788290895041002e-09
Rbbr52 netL52 0 102762362.20681782
Cbr52 netL52 0 -1.5906866940850275e-25

* Branch 53
Rabr53 node_4 netRa53 1695324.6549984263
Lbr53 netRa53 netL53 5.863768135086807e-10
Rbbr53 netL53 0 -1847517.4394696865
Cbr53 netL53 0 1.8753422013660816e-22

* Branch 54
Rabr54 node_4 netRa54 5461.280213636629
Lbr54 netRa54 netL54 1.612187356373453e-11
Rbbr54 netL54 0 -82341.66368616356
Cbr54 netL54 0 3.635460653173374e-20

* Branch 55
Rabr55 node_4 netRa55 -4004.1673948390544
Lbr55 netRa55 netL55 -6.145621583073731e-11
Rbbr55 netL55 0 776670.1395070328
Cbr55 netL55 0 -2.1144423788245996e-20

* Branch 56
Rabr56 node_4 netRa56 -17380.75666836499
Lbr56 netRa56 netL56 1.815437027384519e-11
Rbbr56 netL56 0 55576.32535957208
Cbr56 netL56 0 1.8711444722308947e-20

* Branch 57
Rabr57 node_4 netRa57 8647.8991292653
Lbr57 netRa57 netL57 8.999529603083202e-12
Rbbr57 netL57 0 -40453.78246976715
Cbr57 netL57 0 2.5831315726264915e-20

* Branch 58
Rabr58 node_4 netRa58 -60950.99602823883
Lbr58 netRa58 netL58 7.337961100099238e-11
Rbbr58 netL58 0 282413.49627232435
Cbr58 netL58 0 4.24378433741014e-21

* Branch 59
Rabr59 node_4 netRa59 191574.34176365272
Lbr59 netRa59 netL59 -4.8337638151908764e-11
Rbbr59 netL59 0 -209701.17146870572
Cbr59 netL59 0 -1.202103134783471e-21

* Branch 60
Rabr60 node_4 netRa60 -734342.028839768
Lbr60 netRa60 netL60 -3.159086288324114e-10
Rbbr60 netL60 0 1019771.8030200866
Cbr60 netL60 0 -4.225095539090079e-22

* Branch 61
Rabr61 node_4 netRa61 172780.9834070307
Lbr61 netRa61 netL61 -4.442899272794209e-11
Rbbr61 netL61 0 -205873.95157605878
Cbr61 netL61 0 -1.2478914712995809e-21

* Branch 62
Rabr62 node_4 netRa62 -17217.657173000447
Lbr62 netRa62 netL62 -9.639219171550045e-11
Rbbr62 netL62 0 319765.4394755463
Cbr62 netL62 0 -1.784842338813975e-20

* Branch 63
Rabr63 node_4 netRa63 -126124.06397684096
Lbr63 netRa63 netL63 -1.3379412286131487e-10
Rbbr63 netL63 0 201593.63227523008
Cbr63 netL63 0 -5.2811840412370504e-21

* Branch 64
Rabr64 node_4 netRa64 12850.041294104938
Lbr64 netRa64 netL64 -5.0867653389105505e-11
Rbbr64 netL64 0 -99457.29715423589
Cbr64 netL64 0 -3.931173644695974e-20

* Branch 65
Rabr65 node_4 netRa65 1797131.1273758477
Lbr65 netRa65 netL65 -3.1527533090491626e-10
Rbbr65 netL65 0 -1853581.7432960507
Cbr65 netL65 0 -9.459521196098798e-23

* Branch 66
Rabr66 node_4 netRa66 7710.074467511047
Lbr66 netRa66 netL66 -5.1296798832871596e-11
Rbbr66 netL66 0 -147566.73324587863
Cbr66 netL66 0 -4.420199720751231e-20

* Branch 67
Rabr67 node_4 netRa67 -2844549.541301588
Lbr67 netRa67 netL67 -3.4691086586554274e-10
Rbbr67 netL67 0 2919693.6319743153
Cbr67 netL67 0 -4.178447902232352e-23

* Branch 68
Rabr68 node_4 netRa68 -10704.938101469623
Lbr68 netRa68 netL68 -1.1455300092058823e-10
Rbbr68 netL68 0 806460.0122709593
Cbr68 netL68 0 -1.3669724109062994e-20

* Branch 69
Rabr69 node_4 netRa69 4067.094565674813
Lbr69 netRa69 netL69 -5.416967774959668e-11
Rbbr69 netL69 0 -282859.6126843252
Cbr69 netL69 0 -4.543348963319234e-20

* Branch 70
Rabr70 node_4 netRa70 4407.6553522568865
Lbr70 netRa70 netL70 -3.51074315716726e-11
Rbbr70 netL70 0 -128320.36278356207
Cbr70 netL70 0 -6.079075762048101e-20

* Branch 71
Rabr71 node_4 netRa71 528361.1633640461
Lbr71 netRa71 netL71 -1.0427688316109261e-10
Rbbr71 netL71 0 -591215.0890491639
Cbr71 netL71 0 -3.3366032535934136e-22

* Branch 72
Rabr72 node_4 netRa72 1240.2217457560855
Lbr72 netRa72 netL72 8.61758179145703e-12
Rbbr72 netL72 0 -31497.01508192258
Cbr72 netL72 0 2.2381880189202383e-19

* Branch 73
Rabr73 node_4 netRa73 3492.8209914900144
Lbr73 netRa73 netL73 1.0475244007685773e-11
Rbbr73 netL73 0 -72514.8166297562
Cbr73 netL73 0 4.155947465783132e-20

* Branch 74
Rabr74 node_4 netRa74 61665.196863323275
Lbr74 netRa74 netL74 3.804024006393312e-11
Rbbr74 netL74 0 -99991.94933840747
Cbr74 netL74 0 6.1748144642763096e-21

* Branch 75
Rabr75 node_4 netRa75 101.06683740979217
Lbr75 netRa75 netL75 2.495543370008139e-12
Rbbr75 netL75 0 -77875.17585242329
Cbr75 netL75 0 3.262990037672225e-19

* Branch 76
Rabr76 node_4 netRa76 79645.00886579951
Lbr76 netRa76 netL76 -5.993038823630417e-11
Rbbr76 netL76 0 -121270.42271469039
Cbr76 netL76 0 -6.199678048767445e-21

* Branch 77
Rabr77 node_4 netRa77 11659.894519892014
Lbr77 netRa77 netL77 2.0920976940453348e-11
Rbbr77 netL77 0 -74756.17153646189
Cbr77 netL77 0 2.4036876112774656e-20

* Branch 78
Rabr78 node_4 netRa78 109988.27500281889
Lbr78 netRa78 netL78 -8.409992998579909e-11
Rbbr78 netL78 0 -170610.13562465706
Cbr78 netL78 0 -4.479341314470999e-21

* Branch 79
Rabr79 node_4 netRa79 -120153.1657694788
Lbr79 netRa79 netL79 -1.6396249402809245e-10
Rbbr79 netL79 0 247241.12653845715
Cbr79 netL79 0 -5.523847417431434e-21

* Branch 80
Rabr80 node_4 netRa80 468907.27826552076
Lbr80 netRa80 netL80 -1.8830996787269248e-10
Rbbr80 netL80 0 -715174.6620083784
Cbr80 netL80 0 -5.613984798092325e-22

* Branch 81
Rabr81 node_4 netRa81 163331.33602774082
Lbr81 netRa81 netL81 5.48049546905956e-10
Rbbr81 netL81 0 -2989843.3975109565
Cbr81 netL81 0 1.1242990732979733e-21

* Branch 82
Rabr82 node_4 netRa82 -97230.7296125923
Lbr82 netRa82 netL82 -9.45686589405192e-11
Rbbr82 netL82 0 153168.35878270635
Cbr82 netL82 0 -6.350125963529831e-21

* Branch 83
Rabr83 node_4 netRa83 508991.6027370803
Lbr83 netRa83 netL83 1.462651345332198e-10
Rbbr83 netL83 0 -620059.9342945096
Cbr83 netL83 0 4.63452502328521e-22

* Branch 84
Rabr84 node_4 netRa84 -12436.77686620215
Lbr84 netRa84 netL84 -2.5240614374872512e-11
Rbbr84 netL84 0 38285.08937662368
Cbr84 netL84 0 -5.301910855355916e-20

* Branch 85
Rabr85 node_4 netRa85 -114393.58138192171
Lbr85 netRa85 netL85 -1.081638007955207e-10
Rbbr85 netL85 0 174509.90137390522
Cbr85 netL85 0 -5.418836716994665e-21

* Branch 86
Rabr86 node_4 netRa86 48408.60246239056
Lbr86 netRa86 netL86 -8.706402348946678e-11
Rbbr86 netL86 0 -550324.8704928635
Cbr86 netL86 0 -3.2663825484439827e-21

* Branch 87
Rabr87 node_4 netRa87 -169196.50826332482
Lbr87 netRa87 netL87 4.0547424537622864e-11
Rbbr87 netL87 0 199905.52953725637
Cbr87 netL87 0 1.1987017489690974e-21

* Branch 88
Rabr88 node_4 netRa88 27744.31492902792
Lbr88 netRa88 netL88 -4.941489725597637e-11
Rbbr88 netL88 0 -192969.1432689673
Cbr88 netL88 0 -9.219065071399487e-21

* Branch 89
Rabr89 node_4 netRa89 -53972010.21073223
Lbr89 netRa89 netL89 1.4940852392601807e-09
Rbbr89 netL89 0 54096389.31253656
Cbr89 netL89 0 5.117095582034362e-25

* Branch 90
Rabr90 node_4 netRa90 -7558.644237948751
Lbr90 netRa90 netL90 3.0711799545324636e-11
Rbbr90 netL90 0 201523.81678729423
Cbr90 netL90 0 2.0051549826502627e-20

* Branch 91
Rabr91 node_4 netRa91 138478.98910811412
Lbr91 netRa91 netL91 8.559266563815964e-11
Rbbr91 netL91 0 -194082.32546632513
Cbr91 netL91 0 3.1877735336142205e-21

* Branch 92
Rabr92 node_4 netRa92 1309256.4156175666
Lbr92 netRa92 netL92 1.2575052743594022e-10
Rbbr92 netL92 0 -1339121.4021675007
Cbr92 netL92 0 7.174153378148997e-23

* Branch 93
Rabr93 node_4 netRa93 -14881.840096678172
Lbr93 netRa93 netL93 -9.353791049547533e-12
Rbbr93 netL93 0 34836.38339736622
Cbr93 netL93 0 -1.80789275645143e-20

* Branch 94
Rabr94 node_4 netRa94 -1708688.094583471
Lbr94 netRa94 netL94 -2.358910719192249e-10
Rbbr94 netL94 0 1724612.9529221295
Cbr94 netL94 0 -8.009144294143196e-23

* Branch 95
Rabr95 node_4 netRa95 -315653.58240521426
Lbr95 netRa95 netL95 -7.978970039312194e-11
Rbbr95 netL95 0 387117.103407958
Cbr95 netL95 0 -6.536548632402539e-22

* Branch 96
Rabr96 node_4 netRa96 111.83445657902405
Lbr96 netRa96 netL96 1.908882610878602e-13
Rbbr96 netL96 0 -859.4382528685247
Cbr96 netL96 0 2.0199012890885583e-18

* Branch 97
Rabr97 node_4 netRa97 601.5461341208995
Lbr97 netRa97 netL97 7.440151596927572e-14
Rbbr97 netL97 0 -627.1625369767133
Cbr97 netL97 0 1.9763721924589551e-19

* Branch 98
Rabr98 node_4 netRa98 263.30292155507766
Lbr98 netRa98 netL98 6.47631599953394e-14
Rbbr98 netL98 0 -295.06456820498795
Cbr98 netL98 0 8.372944718039989e-19

* Branch 99
Rabr99 node_4 netRa99 -72.94425170999612
Lbr99 netRa99 netL99 1.9886780892324936e-14
Rbbr99 netL99 0 79.62067182288104
Cbr99 netL99 0 3.3071379509486908e-18

.ends


.end
